`timescale 1 ns / 1 ps

module ml_model_stage1 (
    input [286:0] model_inp,
    output [94:0] model_out
);

    // verilator lint_off UNUSEDSIGNAL
    // Explicit quantization operation will drop bits if exists

    wire [4:0] v0; assign v0[4:0] = model_inp[4:0]; // 10.0
    wire [4:0] v1; assign v1[4:0] = model_inp[9:5]; // 10.0
    wire [6:0] v2; shift_adder #(5, 5, 1, 1, 7, -1, 1) op_2 (v0[4:0], v1[4:0], v2[6:0]); // 11.0
    wire [5:0] v3; assign v3[5:0] = model_inp[15:10]; // 10.0
    wire [4:0] v4; assign v4[4:0] = model_inp[20:16]; // 10.0
    wire [6:0] v5; shift_adder #(6, 5, 1, 1, 7, 1, 0) op_5 (v3[5:0], v4[4:0], v5[6:0]); // 11.0
    wire [4:0] v6; assign v6[4:0] = model_inp[25:21]; // 10.0
    wire [3:0] v7; assign v7[3:0] = model_inp[29:26]; // 10.0
    wire [6:0] v8; shift_adder #(5, 4, 1, 1, 7, -1, 0) op_8 (v6[4:0], v7[3:0], v8[6:0]); // 11.0
    wire [4:0] v9; assign v9[4:0] = model_inp[34:30]; // 10.0
    wire [4:0] v10; assign v10[4:0] = model_inp[39:35]; // 10.0
    wire [5:0] v11; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_11 (v9[4:0], v10[4:0], v11[5:0]); // 11.0
    wire [4:0] v12; assign v12[4:0] = model_inp[44:40]; // 10.0
    wire [4:0] v13; assign v13[4:0] = model_inp[49:45]; // 10.0
    wire [6:0] v14; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_14 (v12[4:0], v13[4:0], v14[6:0]); // 11.0
    wire [4:0] v15; assign v15[4:0] = model_inp[54:50]; // 10.0
    wire [5:0] v16; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_16 (v4[4:0], v15[4:0], v16[5:0]); // 11.0
    wire [5:0] v17; assign v17[5:0] = model_inp[60:55]; // 10.0
    wire [4:0] v18; assign v18[4:0] = model_inp[65:61]; // 10.0
    wire [6:0] v19; shift_adder #(6, 5, 1, 1, 7, -1, 0) op_19 (v17[5:0], v18[4:0], v19[6:0]); // 11.0
    wire [4:0] v20; assign v20[4:0] = model_inp[70:66]; // 10.0
    wire [6:0] v21; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_21 (v12[4:0], v20[4:0], v21[6:0]); // 11.0
    wire [5:0] v22; assign v22[5:0] = model_inp[76:71]; // 10.0
    wire [5:0] v23; assign v23[5:0] = model_inp[82:77]; // 10.0
    wire [7:0] v24; shift_adder #(6, 6, 1, 1, 8, 1, 0) op_24 (v22[5:0], v23[5:0], v24[7:0]); // 11.0
    wire [4:0] v25; assign v25[4:0] = model_inp[87:83]; // 10.0
    wire [5:0] v26; assign v26[5:0] = model_inp[93:88]; // 10.0
    wire [6:0] v27; shift_adder #(5, 6, 1, 1, 7, 0, 0) op_27 (v25[4:0], v26[5:0], v27[6:0]); // 11.0
    wire [4:0] v28; assign v28[4:0] = model_inp[98:94]; // 10.0
    wire [7:0] v29; shift_adder #(5, 5, 1, 1, 8, -2, 1) op_29 (v28[4:0], v4[4:0], v29[7:0]); // 11.0
    wire [8:0] v30; shift_adder #(5, 5, 1, 1, 9, -3, 0) op_30 (v18[4:0], v13[4:0], v30[8:0]); // 11.0
    wire [4:0] v31; assign v31[4:0] = model_inp[103:99]; // 10.0
    wire [5:0] v32; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_32 (v31[4:0], v28[4:0], v32[5:0]); // 11.0
    wire [4:0] v33; assign v33[4:0] = model_inp[108:104]; // 10.0
    wire [4:0] v34; assign v34[4:0] = model_inp[113:109]; // 10.0
    wire [5:0] v35; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_35 (v33[4:0], v34[4:0], v35[5:0]); // 11.0
    wire [6:0] v36; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_36 (v22[5:0], v23[5:0], v36[6:0]); // 11.0
    wire [5:0] v37; assign v37[5:0] = model_inp[119:114]; // 10.0
    wire [5:0] v38; assign v38[5:0] = model_inp[125:120]; // 10.0
    wire [7:0] v39; shift_adder #(6, 6, 1, 1, 8, 1, 0) op_39 (v37[5:0], v38[5:0], v39[7:0]); // 11.0
    wire [4:0] v40; assign v40[4:0] = model_inp[130:126]; // 10.0
    wire [4:0] v41; assign v41[4:0] = model_inp[135:131]; // 10.0
    wire [5:0] v42; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_42 (v40[4:0], v41[4:0], v42[5:0]); // 11.0
    wire [5:0] v43; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_43 (v31[4:0], v28[4:0], v43[5:0]); // 11.0
    wire [4:0] v44; assign v44[4:0] = model_inp[140:136]; // 10.0
    wire [6:0] v45; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_45 (v20[4:0], v44[4:0], v45[6:0]); // 11.0
    wire [7:0] v46; shift_adder #(5, 5, 1, 1, 8, -2, 1) op_46 (v41[4:0], v34[4:0], v46[7:0]); // 11.0
    wire [6:0] v47; shift_adder #(5, 5, 1, 1, 7, -1, 0) op_47 (v33[4:0], v25[4:0], v47[6:0]); // 11.0
    wire [4:0] v48; assign v48[4:0] = model_inp[145:141]; // 10.0
    wire [6:0] v49; shift_adder #(5, 6, 1, 1, 7, 0, 0) op_49 (v48[4:0], v22[5:0], v49[6:0]); // 11.0
    wire [4:0] v50; assign v50[4:0] = model_inp[150:146]; // 10.0
    wire [7:0] v51; shift_adder #(5, 5, 1, 1, 8, -2, 1) op_51 (v50[4:0], v28[4:0], v51[7:0]); // 11.0
    wire [6:0] v52; shift_adder #(5, 5, 1, 1, 7, -1, 0) op_52 (v31[4:0], v44[4:0], v52[6:0]); // 11.0
    wire [6:0] v53; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_53 (v37[5:0], v38[5:0], v53[6:0]); // 11.0
    wire [5:0] v54; assign v54[5:0] = model_inp[156:151]; // 10.0
    wire [5:0] v55; assign v55[5:0] = model_inp[162:157]; // 10.0
    wire [6:0] v56; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_56 (v54[5:0], v55[5:0], v56[6:0]); // 11.0
    wire [4:0] v57; assign v57[4:0] = model_inp[167:163]; // 10.0
    wire [5:0] v58; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_58 (v57[4:0], v50[4:0], v58[5:0]); // 11.0
    wire [5:0] v59; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_59 (v40[4:0], v41[4:0], v59[5:0]); // 11.0
    wire [4:0] v60; assign v60[4:0] = model_inp[172:168]; // 10.0
    wire [2:0] v61; assign v61[2:0] = model_inp[175:173]; // 10.0
    wire [5:0] v62; shift_adder #(5, 3, 1, 0, 6, 1, 1) op_62 (v60[4:0], v61[2:0], v62[5:0]); // 11.0
    wire [5:0] v63; assign v63[5:0] = model_inp[181:176]; // 10.0
    wire [6:0] v64; assign v64[6:0] = model_inp[188:182]; // 10.0
    wire [7:0] v65; shift_adder #(6, 7, 1, 1, 8, -1, 0) op_65 (v63[5:0], v64[6:0], v65[7:0]); // 11.0
    wire [4:0] v66; assign v66[4:0] = model_inp[193:189]; // 10.0
    wire [4:0] v67; assign v67[4:0] = model_inp[198:194]; // 10.0
    wire [6:0] v68; shift_adder #(5, 5, 1, 1, 7, -1, 0) op_68 (v66[4:0], v67[4:0], v68[6:0]); // 11.0
    wire [4:0] v69; assign v69[4:0] = model_inp[203:199]; // 10.0
    wire [4:0] v70; assign v70[4:0] = model_inp[208:204]; // 10.0
    wire [6:0] v71; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_71 (v69[4:0], v70[4:0], v71[6:0]); // 11.0
    wire [5:0] v72; assign v72[5:0] = model_inp[214:209]; // 10.0
    wire [7:0] v73; shift_adder #(5, 6, 1, 1, 8, 1, 0) op_73 (v0[4:0], v72[5:0], v73[7:0]); // 11.0
    wire [5:0] v74; assign v74[5:0] = model_inp[220:215]; // 10.0
    wire [6:0] v75; assign v75[6:0] = model_inp[227:221]; // 10.0
    wire [7:0] v76; shift_adder #(6, 7, 1, 1, 8, 0, 0) op_76 (v74[5:0], v75[6:0], v76[7:0]); // 11.0
    wire [5:0] v77; assign v77[5:0] = model_inp[233:228]; // 10.0
    wire [6:0] v78; shift_adder #(6, 5, 1, 1, 7, 0, 0) op_78 (v77[5:0], v6[4:0], v78[6:0]); // 11.0
    wire [5:0] v79; shift_adder #(5, 3, 1, 0, 6, 1, 1) op_79 (v48[4:0], v61[2:0], v79[5:0]); // 11.0
    wire [7:0] v80; shift_adder #(5, 5, 1, 1, 8, 2, 0) op_80 (v70[4:0], v57[4:0], v80[7:0]); // 11.0
    wire [6:0] v81; assign v81[6:0] = model_inp[240:234]; // 10.0
    wire [7:0] v82; shift_adder #(5, 7, 1, 1, 8, -1, 0) op_82 (v67[4:0], v81[6:0], v82[7:0]); // 11.0
    wire [5:0] v83; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_83 (v60[4:0], v69[4:0], v83[5:0]); // 11.0
    wire [7:0] v84; assign v84[7:0] = model_inp[248:241]; // 10.0
    wire [7:0] v85; shift_adder #(8, 5, 1, 1, 8, 0, 1) op_85 (v84[7:0], v50[4:0], v85[7:0]); // 11.0
    wire [6:0] v86; shift_adder #(6, 5, 1, 1, 7, 1, 0) op_86 (v55[5:0], v66[4:0], v86[6:0]); // 11.0
    wire [6:0] v87; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_87 (v9[4:0], v12[4:0], v87[6:0]); // 11.0
    wire [6:0] v88; shift_adder #(5, 5, 1, 1, 7, -1, 0) op_88 (v13[4:0], v20[4:0], v88[6:0]); // 11.0
    wire [5:0] v89; assign v89[5:0] = model_inp[254:249]; // 10.0
    wire [6:0] v90; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_90 (v89[5:0], v26[5:0], v90[6:0]); // 11.0
    wire [6:0] v91; shift_adder #(5, 4, 1, 1, 7, -1, 1) op_91 (v34[4:0], v7[3:0], v91[6:0]); // 11.0
    wire [6:0] v92; shift_adder #(5, 5, 1, 1, 7, -1, 0) op_92 (v15[4:0], v10[4:0], v92[6:0]); // 11.0
    wire [5:0] v93; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_93 (v33[4:0], v34[4:0], v93[5:0]); // 11.0
    wire [5:0] v94; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_94 (v18[4:0], v4[4:0], v94[5:0]); // 11.0
    wire [6:0] v95; shift_adder #(5, 5, 1, 1, 7, -1, 0) op_95 (v48[4:0], v60[4:0], v95[6:0]); // 11.0
    wire [5:0] v96; assign v96[5:0] = model_inp[260:255]; // 10.0
    wire [6:0] v97; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_97 (v55[5:0], v96[5:0], v97[6:0]); // 11.0
    wire [6:0] v98; shift_adder #(5, 6, 1, 1, 7, -1, 0) op_98 (v69[4:0], v37[5:0], v98[6:0]); // 11.0
    wire [7:0] v99; shift_adder #(5, 5, 1, 1, 8, -2, 1) op_99 (v70[4:0], v41[4:0], v99[7:0]); // 11.0
    wire [6:0] v100; shift_adder #(6, 5, 1, 1, 7, 1, 0) op_100 (v38[5:0], v66[4:0], v100[6:0]); // 11.0
    wire [5:0] v101; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_101 (v70[4:0], v57[4:0], v101[5:0]); // 11.0
    wire [7:0] v102; shift_adder #(5, 5, 1, 1, 8, 2, 0) op_102 (v50[4:0], v40[4:0], v102[7:0]); // 11.0
    wire [6:0] v103; shift_adder #(5, 5, 1, 1, 7, -1, 0) op_103 (v0[4:0], v9[4:0], v103[6:0]); // 11.0
    wire [4:0] v104; assign v104[4:0] = model_inp[265:261]; // 10.0
    wire [5:0] v105; shift_adder #(5, 4, 1, 1, 6, 1, 0) op_105 (v104[4:0], v7[3:0], v105[5:0]); // 11.0
    wire [6:0] v106; assign v106[6:0] = model_inp[272:266]; // 10.0
    wire [7:0] v107; shift_adder #(7, 6, 1, 1, 8, 1, 0) op_107 (v106[6:0], v3[5:0], v107[7:0]); // 11.0
    wire [5:0] v108; shift_adder #(5, 4, 1, 1, 6, 1, 0) op_108 (v6[4:0], v7[3:0], v108[5:0]); // 11.0
    wire [8:0] v109; assign v109[8:0] = model_inp[281:273]; // 10.0
    wire [8:0] v110; shift_adder #(9, 5, 1, 1, 9, 1, 0) op_110 (v109[8:0], v15[4:0], v110[8:0]); // 11.0
    wire [9:0] v111; shift_adder #(7, 7, 1, 1, 10, 2, 0) op_111 (v2[6:0], v5[6:0], v111[9:0]); // 12.0
    wire [7:0] v112; shift_adder #(6, 7, 1, 1, 8, -1, 0) op_112 (v11[5:0], v14[6:0], v112[7:0]); // 12.0
    wire [7:0] v113; shift_adder #(6, 7, 1, 1, 8, 0, 0) op_113 (v16[5:0], v19[6:0], v113[7:0]); // 12.0
    wire [8:0] v114; shift_adder #(7, 8, 1, 1, 9, 0, 0) op_114 (v21[6:0], v24[7:0], v114[8:0]); // 12.0
    wire [7:0] v115; shift_adder #(7, 6, 1, 1, 8, 0, 1) op_115 (v27[6:0], v89[5:0], v115[7:0]); // 12.0
    wire [9:0] v116; shift_adder #(8, 9, 1, 1, 10, -1, 1) op_116 (v29[7:0], v30[8:0], v116[9:0]); // 12.0
    wire [6:0] v117; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_117 (v32[5:0], v35[5:0], v117[6:0]); // 12.0
    wire [8:0] v118; shift_adder #(7, 8, 1, 1, 9, -1, 0) op_118 (v36[6:0], v39[7:0], v118[8:0]); // 12.0
    wire [6:0] v119; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_119 (v42[5:0], v43[5:0], v119[6:0]); // 12.0
    wire [7:0] v120; shift_adder #(7, 6, 1, 1, 8, -1, 1) op_120 (v45[6:0], v26[5:0], v120[7:0]); // 12.0
    wire [8:0] v121; shift_adder #(8, 7, 1, 1, 9, 1, 1) op_121 (v46[7:0], v47[6:0], v121[8:0]); // 12.0
    wire [7:0] v122; shift_adder #(7, 6, 1, 1, 8, -1, 1) op_122 (v49[6:0], v23[5:0], v122[7:0]); // 12.0
    wire [8:0] v123; shift_adder #(8, 7, 1, 1, 9, 1, 1) op_123 (v51[7:0], v52[6:0], v123[8:0]); // 12.0
    wire [7:0] v124; shift_adder #(7, 7, 1, 1, 8, 0, 0) op_124 (v53[6:0], v56[6:0], v124[7:0]); // 12.0
    wire [6:0] v125; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_125 (v58[5:0], v59[5:0], v125[6:0]); // 12.0
    wire [8:0] v126; shift_adder #(6, 8, 1, 1, 9, 0, 0) op_126 (v62[5:0], v65[7:0], v126[8:0]); // 12.0
    wire [8:0] v127; shift_adder #(7, 7, 1, 1, 9, -2, 0) op_127 (v68[6:0], v71[6:0], v127[8:0]); // 12.0
    wire [8:0] v128; shift_adder #(8, 8, 1, 1, 9, 1, 0) op_128 (v73[7:0], v76[7:0], v128[8:0]); // 12.0
    wire [7:0] v129; shift_adder #(6, 6, 1, 1, 8, 1, 1) op_129 (v79[5:0], v96[5:0], v129[7:0]); // 12.0
    wire [8:0] v130; shift_adder #(8, 6, 1, 1, 9, 1, 0) op_130 (v82[7:0], v83[5:0], v130[8:0]); // 12.0
    wire [8:0] v131; shift_adder #(8, 7, 1, 1, 9, -1, 1) op_131 (v85[7:0], v86[6:0], v131[8:0]); // 12.0
    wire [7:0] v132; shift_adder #(7, 6, 1, 1, 8, -1, 1) op_132 (v87[6:0], v3[5:0], v132[7:0]); // 12.0
    wire [8:0] v133; shift_adder #(7, 7, 1, 1, 9, 1, 0) op_133 (v88[6:0], v90[6:0], v133[8:0]); // 12.0
    wire [7:0] v134; shift_adder #(7, 7, 1, 1, 8, 0, 1) op_134 (v91[6:0], v92[6:0], v134[7:0]); // 12.0
    wire [6:0] v135; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_135 (v93[5:0], v94[5:0], v135[6:0]); // 12.0
    wire [8:0] v136; shift_adder #(7, 7, 1, 1, 9, 1, 0) op_136 (v95[6:0], v97[6:0], v136[8:0]); // 12.0
    wire [7:0] v137; shift_adder #(7, 6, 1, 1, 8, 1, 1) op_137 (v98[6:0], v54[5:0], v137[7:0]); // 12.0
    wire [8:0] v138; shift_adder #(8, 7, 1, 1, 9, -1, 1) op_138 (v99[7:0], v100[6:0], v138[8:0]); // 12.0
    wire [7:0] v139; shift_adder #(6, 8, 1, 1, 8, 0, 0) op_139 (v101[5:0], v102[7:0], v139[7:0]); // 12.0
    wire [4:0] v140; assign v140[4:0] = model_inp[286:282]; // 10.0
    wire [7:0] v141; shift_adder #(7, 5, 1, 1, 8, 1, 1) op_141 (v103[6:0], v140[4:0], v141[7:0]); // 12.0
    wire [8:0] v142; shift_adder #(6, 8, 1, 1, 9, -2, 0) op_142 (v105[5:0], v107[7:0], v142[8:0]); // 12.0
    wire [8:0] v143; shift_adder #(6, 9, 1, 1, 9, -1, 0) op_143 (v108[5:0], v110[8:0], v143[8:0]); // 12.0
    wire [9:0] v144; shift_adder #(10, 7, 1, 1, 10, 2, 1) op_144 (v111[9:0], v8[6:0], v144[9:0]); // 13.0
    wire [8:0] v145; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_145 (v112[7:0], v113[7:0], v145[8:0]); // 13.0
    wire [9:0] v146; shift_adder #(9, 8, 1, 1, 10, 1, 0) op_146 (v114[8:0], v115[7:0], v146[9:0]); // 13.0
    wire [9:0] v147; shift_adder #(10, 7, 1, 1, 10, 1, 1) op_147 (v116[9:0], v117[6:0], v147[9:0]); // 13.0
    wire [9:0] v148; shift_adder #(9, 7, 1, 1, 10, 0, 1) op_148 (v118[8:0], v119[6:0], v148[9:0]); // 13.0
    wire [9:0] v149; shift_adder #(8, 9, 1, 1, 10, 1, 0) op_149 (v120[7:0], v121[8:0], v149[9:0]); // 13.0
    wire [9:0] v150; shift_adder #(8, 9, 1, 1, 10, 1, 0) op_150 (v122[7:0], v123[8:0], v150[9:0]); // 13.0
    wire [9:0] v151; shift_adder #(8, 7, 1, 1, 10, -1, 1) op_151 (v124[7:0], v125[6:0], v151[9:0]); // 13.0
    wire [9:0] v152; shift_adder #(9, 9, 1, 1, 10, -1, 1) op_152 (v126[8:0], v127[8:0], v152[9:0]); // 13.0
    wire [9:0] v153; shift_adder #(10, 3, 1, 0, 10, 0, 1) op_153 (v152[9:0], 3'b101, v153[9:0]); // 13.0
    wire [8:0] v154; assign v154[8:0] = v153[8:0] & {9{~v153[9]}}; // 13.0
    wire [8:0] v155; shift_adder #(9, 4, 0, 0, 9, 0, 0) op_155 (v154[8:0], 4'b1000, v155[8:0]); // 13.0
    wire [3:0] v156; assign v156[3:0] = v155[7:4]; // 13.0
    wire [9:0] v157; shift_adder #(9, 7, 1, 1, 10, 0, 1) op_157 (v128[8:0], v78[6:0], v157[9:0]); // 13.0
    wire [10:0] v158; shift_adder #(10, 3, 1, 0, 11, -1, 1) op_158 (v157[9:0], 3'b101, v158[10:0]); // 13.0
    wire [8:0] v159; assign v159[8:0] = v158[8:0] & {9{~v158[10]}}; // 13.0
    wire [8:0] v160; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_160 (v159[8:0], 3'b100, v160[8:0]); // 13.0
    wire [5:0] v161; assign v161[5:0] = v160[8:3]; // 13.0
    wire [8:0] v162; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_162 (v129[7:0], v80[7:0], v162[8:0]); // 13.0
    wire [10:0] v163; shift_adder #(9, 9, 1, 1, 11, -1, 0) op_163 (v130[8:0], v131[8:0], v163[10:0]); // 13.0
    wire [9:0] v164; shift_adder #(8, 9, 1, 1, 10, 1, 0) op_164 (v132[7:0], v133[8:0], v164[9:0]); // 13.0
    wire [8:0] v165; shift_adder #(8, 7, 1, 1, 9, -1, 1) op_165 (v134[7:0], v135[6:0], v165[8:0]); // 13.0
    wire [9:0] v166; shift_adder #(9, 8, 1, 1, 10, 0, 0) op_166 (v136[8:0], v137[7:0], v166[9:0]); // 13.0
    wire [9:0] v167; shift_adder #(9, 8, 1, 1, 10, 1, 1) op_167 (v138[8:0], v139[7:0], v167[9:0]); // 13.0
    wire [9:0] v168; shift_adder #(8, 9, 1, 1, 10, 0, 0) op_168 (v141[7:0], v142[8:0], v168[9:0]); // 13.0
    wire [10:0] v169; shift_adder #(10, 9, 1, 1, 11, 1, 0) op_169 (v144[9:0], v145[8:0], v169[10:0]); // 14.0
    wire [10:0] v170; shift_adder #(11, 3, 1, 0, 11, 0, 1) op_170 (v169[10:0], 3'b101, v170[10:0]); // 14.0
    wire [9:0] v171; assign v171[9:0] = v170[9:0] & {10{~v170[10]}}; // 14.0
    wire [9:0] v172; shift_adder #(10, 3, 0, 0, 10, 0, 0) op_172 (v171[9:0], 3'b100, v172[9:0]); // 14.0
    wire [5:0] v173; assign v173[5:0] = v172[8:3]; // 14.0
    wire [10:0] v174; shift_adder #(10, 10, 1, 1, 11, -1, 0) op_174 (v146[9:0], v147[9:0], v174[10:0]); // 14.0
    wire [10:0] v175; shift_adder #(11, 3, 1, 0, 11, 0, 1) op_175 (v174[10:0], 3'b101, v175[10:0]); // 14.0
    wire [9:0] v176; assign v176[9:0] = v175[9:0] & {10{~v175[10]}}; // 14.0
    wire [9:0] v177; shift_adder #(10, 3, 0, 0, 10, 0, 0) op_177 (v176[9:0], 3'b100, v177[9:0]); // 14.0
    wire [5:0] v178; assign v178[5:0] = v177[8:3]; // 14.0
    wire [11:0] v179; shift_adder #(10, 10, 1, 1, 12, -1, 0) op_179 (v148[9:0], v149[9:0], v179[11:0]); // 14.0
    wire [11:0] v180; shift_adder #(12, 3, 1, 0, 12, 0, 1) op_180 (v179[11:0], 3'b101, v180[11:0]); // 14.0
    wire [9:0] v181; assign v181[9:0] = v180[9:0] & {10{~v180[11]}}; // 14.0
    wire [10:0] v182; shift_adder #(10, 3, 0, 0, 11, 0, 0) op_182 (v181[9:0], 3'b100, v182[10:0]); // 14.0
    wire [5:0] v183; assign v183[5:0] = v182[8:3]; // 14.0
    wire [11:0] v184; shift_adder #(10, 10, 1, 1, 12, 1, 0) op_184 (v150[9:0], v151[9:0], v184[11:0]); // 14.0
    wire [11:0] v185; shift_adder #(12, 3, 1, 0, 12, 0, 1) op_185 (v184[11:0], 3'b101, v185[11:0]); // 14.0
    wire [10:0] v186; assign v186[10:0] = v185[10:0] & {11{~v185[11]}}; // 14.0
    wire [10:0] v187; shift_adder #(11, 3, 0, 0, 11, 0, 0) op_187 (v186[10:0], 3'b100, v187[10:0]); // 14.0
    wire [5:0] v188; assign v188[5:0] = v187[8:3]; // 14.0
    wire [7:0] v189; shift_adder #(4, 6, 1, 1, 8, -3, 0) op_189 (v156[3:0], v161[5:0], v189[7:0]); // 14.0
    wire [10:0] v190; shift_adder #(9, 11, 1, 1, 11, -1, 0) op_190 (v162[8:0], v163[10:0], v190[10:0]); // 14.0
    wire [10:0] v191; shift_adder #(11, 3, 1, 0, 11, 0, 1) op_191 (v190[10:0], 3'b101, v191[10:0]); // 14.0
    wire [9:0] v192; assign v192[9:0] = v191[9:0] & {10{~v191[10]}}; // 14.0
    wire [9:0] v193; shift_adder #(10, 3, 0, 0, 10, 0, 0) op_193 (v192[9:0], 3'b100, v193[9:0]); // 14.0
    wire [5:0] v194; assign v194[5:0] = v193[8:3]; // 14.0
    wire [10:0] v195; shift_adder #(10, 9, 1, 1, 11, 1, 0) op_195 (v164[9:0], v165[8:0], v195[10:0]); // 14.0
    wire [10:0] v196; shift_adder #(11, 3, 1, 0, 11, 0, 1) op_196 (v195[10:0], 3'b101, v196[10:0]); // 14.0
    wire [9:0] v197; assign v197[9:0] = v196[9:0] & {10{~v196[10]}}; // 14.0
    wire [9:0] v198; shift_adder #(10, 3, 0, 0, 10, 0, 0) op_198 (v197[9:0], 3'b100, v198[9:0]); // 14.0
    wire [5:0] v199; assign v199[5:0] = v198[8:3]; // 14.0
    wire [11:0] v200; shift_adder #(10, 10, 1, 1, 12, -1, 0) op_200 (v166[9:0], v167[9:0], v200[11:0]); // 14.0
    wire [11:0] v201; shift_adder #(12, 3, 1, 0, 12, 0, 1) op_201 (v200[11:0], 3'b101, v201[11:0]); // 14.0
    wire [9:0] v202; assign v202[9:0] = v201[9:0] & {10{~v201[11]}}; // 14.0
    wire [10:0] v203; shift_adder #(10, 3, 0, 0, 11, 0, 0) op_203 (v202[9:0], 3'b100, v203[10:0]); // 14.0
    wire [5:0] v204; assign v204[5:0] = v203[8:3]; // 14.0
    wire [10:0] v205; shift_adder #(10, 9, 1, 1, 11, -1, 1) op_205 (v168[9:0], v143[8:0], v205[10:0]); // 14.0
    wire [10:0] v206; shift_adder #(11, 3, 1, 0, 11, 0, 1) op_206 (v205[10:0], 3'b101, v206[10:0]); // 14.0
    wire [9:0] v207; assign v207[9:0] = v206[9:0] & {10{~v206[10]}}; // 14.0
    wire [9:0] v208; shift_adder #(10, 3, 0, 0, 10, 0, 0) op_208 (v207[9:0], 3'b100, v208[9:0]); // 14.0
    wire [5:0] v209; assign v209[5:0] = v208[8:3]; // 14.0
    wire [7:0] v210; shift_adder #(6, 6, 1, 1, 8, -1, 0) op_210 (v173[5:0], v178[5:0], v210[7:0]); // 15.0
    wire [7:0] v211; shift_adder #(6, 6, 1, 1, 8, 1, 1) op_211 (v183[5:0], v188[5:0], v211[7:0]); // 15.0
    wire [6:0] v212; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_212 (v199[5:0], v183[5:0], v212[6:0]); // 15.0
    wire [6:0] v213; shift_adder #(6, 4, 1, 1, 7, 2, 1) op_213 (v204[5:0], v156[3:0], v213[6:0]); // 15.0
    wire [7:0] v214; shift_adder #(6, 6, 1, 1, 8, 1, 1) op_214 (v161[5:0], v194[5:0], v214[7:0]); // 15.0
    wire [6:0] v215; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_215 (v178[5:0], v188[5:0], v215[6:0]); // 15.0
    wire [6:0] v216; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_216 (v161[5:0], v194[5:0], v216[6:0]); // 15.0
    wire [8:0] v217; shift_adder #(6, 6, 1, 1, 9, -2, 1) op_217 (v209[5:0], v209[5:0], v217[8:0]); // 15.0
    wire [6:0] v218; shift_adder #(6, 6, 1, 1, 7, 0, 1) op_218 (v173[5:0], v204[5:0], v218[6:0]); // 15.0
    wire [6:0] v219; shift_adder #(6, 4, 1, 1, 7, 1, 0) op_219 (v183[5:0], v156[3:0], v219[6:0]); // 15.0
    wire [6:0] v220; shift_adder #(6, 4, 1, 1, 7, 1, 0) op_220 (v173[5:0], v156[3:0], v220[6:0]); // 15.0
    wire [7:0] v221; shift_adder #(6, 6, 1, 1, 8, 1, 1) op_221 (v194[5:0], v161[5:0], v221[7:0]); // 15.0
    wire [6:0] v222; shift_adder #(6, 4, 1, 1, 7, 2, 1) op_222 (v178[5:0], v156[3:0], v222[6:0]); // 15.0
    wire [7:0] v223; shift_adder #(6, 6, 1, 1, 8, 1, 0) op_223 (v188[5:0], v183[5:0], v223[7:0]); // 15.0
    wire [6:0] v224; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_224 (v209[5:0], v199[5:0], v224[6:0]); // 15.0
    wire [8:0] v225; shift_adder #(6, 6, 1, 1, 9, -2, 1) op_225 (v194[5:0], v161[5:0], v225[8:0]); // 15.0
    wire [7:0] v226; shift_adder #(6, 6, 1, 1, 8, -1, 1) op_226 (v194[5:0], v178[5:0], v226[7:0]); // 15.0
    wire [8:0] v227; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_227 (v211[7:0], v189[7:0], v227[8:0]); // 16.0
    wire [7:0] v228; shift_adder #(6, 7, 1, 1, 8, 0, 1) op_228 (v194[5:0], v212[6:0], v228[7:0]); // 16.0
    wire [8:0] v229; shift_adder #(7, 8, 1, 1, 9, 1, 0) op_229 (v213[6:0], v214[7:0], v229[8:0]); // 16.0
    wire [8:0] v230; shift_adder #(7, 6, 1, 1, 9, 2, 1) op_230 (v216[6:0], v161[5:0], v230[8:0]); // 16.0
    wire [8:0] v231; shift_adder #(4, 9, 1, 1, 9, -2, 0) op_231 (v156[3:0], v217[8:0], v231[8:0]); // 16.0
    wire [8:0] v232; shift_adder #(6, 7, 1, 1, 9, -2, 1) op_232 (v173[5:0], v218[6:0], v232[8:0]); // 16.0
    wire [7:0] v233; shift_adder #(6, 7, 1, 1, 8, -1, 0) op_233 (v199[5:0], v215[6:0], v233[7:0]); // 16.0
    wire [8:0] v234; shift_adder #(7, 7, 1, 1, 9, -2, 1) op_234 (v219[6:0], v220[6:0], v234[8:0]); // 16.0
    wire [7:0] v235; shift_adder #(8, 6, 1, 1, 8, 0, 1) op_235 (v221[7:0], v209[5:0], v235[7:0]); // 16.0
    wire [8:0] v236; shift_adder #(7, 8, 1, 1, 9, 1, 0) op_236 (v222[6:0], v223[7:0], v236[8:0]); // 16.0
    wire [8:0] v237; shift_adder #(7, 8, 1, 1, 9, -1, 0) op_237 (v218[6:0], v214[7:0], v237[8:0]); // 16.0
    wire [9:0] v238; shift_adder #(9, 7, 1, 1, 10, 1, 0) op_238 (v217[8:0], v222[6:0], v238[9:0]); // 16.0
    wire [8:0] v239; shift_adder #(7, 7, 1, 1, 9, 1, 1) op_239 (v218[6:0], v215[6:0], v239[8:0]); // 16.0
    wire [7:0] v240; shift_adder #(7, 7, 1, 1, 8, 0, 0) op_240 (v216[6:0], v219[6:0], v240[7:0]); // 16.0
    wire [8:0] v241; shift_adder #(9, 8, 1, 1, 9, 0, 1) op_241 (v225[8:0], v210[7:0], v241[8:0]); // 16.0
    wire [7:0] v242; shift_adder #(6, 7, 1, 1, 8, 0, 1) op_242 (v161[5:0], v219[6:0], v242[7:0]); // 16.0
    wire [7:0] v243; shift_adder #(6, 7, 1, 1, 8, 0, 0) op_243 (v194[5:0], v224[6:0], v243[7:0]); // 16.0
    wire [7:0] v244; shift_adder #(6, 8, 1, 1, 8, 0, 0) op_244 (v183[5:0], v214[7:0], v244[7:0]); // 16.0
    wire [7:0] v245; shift_adder #(8, 6, 1, 1, 8, 0, 1) op_245 (v226[7:0], v204[5:0], v245[7:0]); // 16.0
    wire [9:0] v246; shift_adder #(8, 9, 1, 1, 10, -1, 0) op_246 (v210[7:0], v227[8:0], v246[9:0]); // 17.0
    wire [8:0] v247; shift_adder #(8, 7, 1, 1, 9, 1, 1) op_247 (v228[7:0], v215[6:0], v247[8:0]); // 17.0
    wire [9:0] v248; shift_adder #(9, 9, 1, 1, 10, 0, 1) op_248 (v230[8:0], v231[8:0], v248[9:0]); // 17.0
    wire [9:0] v249; shift_adder #(9, 8, 1, 1, 10, 0, 0) op_249 (v232[8:0], v233[7:0], v249[9:0]); // 17.0
    wire [8:0] v250; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_250 (v235[7:0], v233[7:0], v250[8:0]); // 17.0
    wire [10:0] v251; shift_adder #(9, 9, 1, 1, 11, 1, 1) op_251 (v236[8:0], v237[8:0], v251[10:0]); // 17.0
    wire [9:0] v252; shift_adder #(9, 7, 1, 1, 10, 1, 1) op_252 (v239[8:0], v224[6:0], v252[9:0]); // 17.0
    wire [9:0] v253; shift_adder #(9, 9, 1, 1, 10, 0, 1) op_253 (v241[8:0], v231[8:0], v253[9:0]); // 17.0
    wire [10:0] v254; shift_adder #(10, 5, 1, 0, 11, -1, 0) op_254 (v253[9:0], 5'b10001, v254[10:0]); // 17.0
    wire [5:0] v255; assign v255[5:0] = v254[8:3]; // 17.0
    wire [8:0] v256; shift_adder #(8, 8, 1, 1, 9, -1, 1) op_256 (v242[7:0], v243[7:0], v256[8:0]); // 17.0
    wire [8:0] v257; shift_adder #(7, 8, 1, 1, 9, 0, 0) op_257 (v224[6:0], v244[7:0], v257[8:0]); // 17.0
    wire [8:0] v258; shift_adder #(8, 7, 1, 1, 9, 0, 1) op_258 (v245[7:0], v220[6:0], v258[8:0]); // 17.0
    wire [10:0] v259; shift_adder #(10, 8, 1, 1, 11, 2, 1) op_259 (v246[9:0], v228[7:0], v259[10:0]); // 18.0
    wire [5:0] v260; assign v260[5:0] = v259[8:3]; // 18.0
    wire [9:0] v261; shift_adder #(9, 9, 1, 1, 10, 0, 0) op_261 (v229[8:0], v247[8:0], v261[9:0]); // 18.0
    wire [9:0] v262; shift_adder #(10, 4, 1, 0, 10, 0, 0) op_262 (v261[9:0], 4'b1110, v262[9:0]); // 18.0
    wire [5:0] v263; assign v263[5:0] = v262[7:2]; // 18.0
    wire [10:0] v264; shift_adder #(10, 10, 1, 1, 11, 0, 1) op_264 (v248[9:0], v249[9:0], v264[10:0]); // 18.0
    wire [10:0] v265; shift_adder #(11, 2, 1, 0, 11, 0, 1) op_265 (v264[10:0], 2'b10, v265[10:0]); // 18.0
    wire [6:0] v266; assign v266[6:0] = v265[8:2]; // 18.0
    wire [9:0] v267; shift_adder #(9, 9, 1, 1, 10, 0, 0) op_267 (v234[8:0], v250[8:0], v267[9:0]); // 18.0
    wire [10:0] v268; shift_adder #(10, 3, 1, 0, 11, -1, 1) op_268 (v267[9:0], 3'b101, v268[10:0]); // 18.0
    wire [6:0] v269; assign v269[6:0] = v268[9:3]; // 18.0
    wire [11:0] v270; shift_adder #(11, 10, 1, 1, 12, 1, 1) op_270 (v251[10:0], v238[9:0], v270[11:0]); // 18.0
    wire [11:0] v271; shift_adder #(12, 4, 1, 0, 12, 0, 0) op_271 (v270[11:0], 4'b1011, v271[11:0]); // 18.0
    wire [5:0] v272; assign v272[5:0] = v271[8:3]; // 18.0
    wire [9:0] v273; shift_adder #(10, 8, 1, 1, 10, 0, 1) op_273 (v252[9:0], v240[7:0], v273[9:0]); // 18.0
    wire [9:0] v274; shift_adder #(10, 2, 1, 0, 10, 0, 1) op_274 (v273[9:0], 2'b11, v274[9:0]); // 18.0
    wire [6:0] v275; assign v275[6:0] = v274[8:2]; // 18.0
    wire [9:0] v276; shift_adder #(9, 9, 1, 1, 10, 0, 1) op_276 (v256[8:0], v232[8:0], v276[9:0]); // 18.0
    wire [10:0] v277; shift_adder #(10, 3, 1, 0, 11, -1, 0) op_277 (v276[9:0], 3'b111, v277[10:0]); // 18.0
    wire [5:0] v278; assign v278[5:0] = v277[8:3]; // 18.0
    wire [9:0] v279; shift_adder #(9, 9, 1, 1, 10, 0, 0) op_279 (v239[8:0], v257[8:0], v279[9:0]); // 18.0
    wire [9:0] v280; shift_adder #(10, 3, 1, 0, 10, 0, 0) op_280 (v279[9:0], 3'b111, v280[9:0]); // 18.0
    wire [5:0] v281; assign v281[5:0] = v280[7:2]; // 18.0
    wire [9:0] v282; shift_adder #(9, 8, 1, 1, 10, -1, 1) op_282 (v258[8:0], v243[7:0], v282[9:0]); // 18.0
    wire [12:0] v283; shift_adder #(10, 5, 1, 0, 13, -3, 0) op_283 (v282[9:0], 5'b11101, v283[12:0]); // 18.0
    wire [5:0] v284; assign v284[5:0] = v283[10:5]; // 18.0
    wire [6:0] v285; shift_adder #(6, 6, 1, 1, 7, 0, 1) op_285 (v260[5:0], v263[5:0], v285[6:0]); // 19.0
    wire [7:0] v286; shift_adder #(7, 7, 1, 1, 8, 0, 1) op_286 (v266[6:0], v269[6:0], v286[7:0]); // 19.0
    wire [7:0] v287; shift_adder #(6, 7, 1, 1, 8, 0, 1) op_287 (v272[5:0], v275[6:0], v287[7:0]); // 19.0
    wire [6:0] v288; shift_adder #(6, 6, 1, 1, 7, 0, 1) op_288 (v255[5:0], v278[5:0], v288[6:0]); // 19.0
    wire [6:0] v289; shift_adder #(6, 6, 1, 1, 7, 0, 1) op_289 (v281[5:0], v284[5:0], v289[6:0]); // 19.0
    wire [5:0] v290; mux #(6, 6, 1, 1, 6, 0, 0) op_290 (v285[6], v263[5:0], v260[5:0], v290[5:0]); // 20.0
    wire [6:0] v291; mux #(7, 7, 1, 1, 7, 0, 0) op_291 (v286[7], v269[6:0], v266[6:0], v291[6:0]); // 20.0
    wire [6:0] v292; mux #(7, 6, 1, 1, 7, 0, 0) op_292 (v287[7], v275[6:0], v272[5:0], v292[6:0]); // 20.0
    wire [5:0] v293; mux #(6, 6, 1, 1, 6, 0, 0) op_293 (v288[6], v278[5:0], v255[5:0], v293[5:0]); // 20.0
    wire [5:0] v294; mux #(6, 6, 1, 1, 6, 0, 0) op_294 (v289[6], v284[5:0], v281[5:0], v294[5:0]); // 20.0

    // verilator lint_on UNUSEDSIGNAL

    assign model_out[5:0] = v290[5:0];
    assign model_out[12:6] = v291[6:0];
    assign model_out[18:13] = v293[5:0];
    assign model_out[24:19] = v294[5:0];
    assign model_out[31:25] = v292[6:0];
    assign model_out[38:32] = v275[6:0];
    assign model_out[45:39] = v269[6:0];
    assign model_out[51:46] = v263[5:0];
    assign model_out[57:52] = v281[5:0];
    assign model_out[63:58] = v255[5:0];
    assign model_out[69:64] = v272[5:0];
    assign model_out[75:70] = v260[5:0];
    assign model_out[81:76] = v284[5:0];
    assign model_out[87:82] = v278[5:0];
    assign model_out[94:88] = v266[6:0];

    endmodule
