`timescale 1 ns / 1 ps

module ml_model_stage0 (
    input [119:0] model_inp,
    output [286:0] model_out
);

    // verilator lint_off UNUSEDSIGNAL
    // Explicit quantization operation will drop bits if exists

    wire [1:0] v0; assign v0[1:0] = model_inp[1:0]; // 0.0
    wire [1:0] v1; assign v1[1:0] = model_inp[3:2]; // 0.0
    wire [1:0] v2; assign v2[1:0] = model_inp[5:4]; // 0.0
    wire [1:0] v3; assign v3[1:0] = model_inp[7:6]; // 0.0
    wire [1:0] v4; assign v4[1:0] = model_inp[9:8]; // 0.0
    wire [1:0] v5; assign v5[1:0] = model_inp[11:10]; // 0.0
    wire [1:0] v6; assign v6[1:0] = model_inp[13:12]; // 0.0
    wire [1:0] v7; assign v7[1:0] = model_inp[15:14]; // 0.0
    wire [1:0] v8; assign v8[1:0] = model_inp[17:16]; // 0.0
    wire [1:0] v9; assign v9[1:0] = model_inp[19:18]; // 0.0
    wire [1:0] v10; assign v10[1:0] = model_inp[21:20]; // 0.0
    wire [1:0] v11; assign v11[1:0] = model_inp[23:22]; // 0.0
    wire [1:0] v12; assign v12[1:0] = model_inp[25:24]; // 0.0
    wire [1:0] v13; assign v13[1:0] = model_inp[27:26]; // 0.0
    wire [1:0] v14; assign v14[1:0] = model_inp[29:28]; // 0.0
    wire [1:0] v15; assign v15[1:0] = model_inp[31:30]; // 0.0
    wire [1:0] v16; assign v16[1:0] = model_inp[33:32]; // 0.0
    wire [1:0] v17; assign v17[1:0] = model_inp[35:34]; // 0.0
    wire [1:0] v18; assign v18[1:0] = model_inp[37:36]; // 0.0
    wire [1:0] v19; assign v19[1:0] = model_inp[39:38]; // 0.0
    wire [1:0] v20; assign v20[1:0] = model_inp[41:40]; // 0.0
    wire [1:0] v21; assign v21[1:0] = model_inp[43:42]; // 0.0
    wire [1:0] v22; assign v22[1:0] = model_inp[45:44]; // 0.0
    wire [1:0] v23; assign v23[1:0] = model_inp[47:46]; // 0.0
    wire [1:0] v24; assign v24[1:0] = model_inp[49:48]; // 0.0
    wire [1:0] v25; assign v25[1:0] = model_inp[51:50]; // 0.0
    wire [1:0] v26; assign v26[1:0] = model_inp[53:52]; // 0.0
    wire [1:0] v27; assign v27[1:0] = model_inp[55:54]; // 0.0
    wire [1:0] v28; assign v28[1:0] = model_inp[57:56]; // 0.0
    wire [1:0] v29; assign v29[1:0] = model_inp[59:58]; // 0.0
    wire [1:0] v30; assign v30[1:0] = model_inp[61:60]; // 0.0
    wire [1:0] v31; assign v31[1:0] = model_inp[63:62]; // 0.0
    wire [1:0] v32; assign v32[1:0] = model_inp[65:64]; // 0.0
    wire [1:0] v33; assign v33[1:0] = model_inp[67:66]; // 0.0
    wire [1:0] v34; assign v34[1:0] = model_inp[69:68]; // 0.0
    wire [1:0] v35; assign v35[1:0] = model_inp[71:70]; // 0.0
    wire [1:0] v36; assign v36[1:0] = model_inp[73:72]; // 0.0
    wire [1:0] v37; assign v37[1:0] = model_inp[75:74]; // 0.0
    wire [1:0] v38; assign v38[1:0] = model_inp[77:76]; // 0.0
    wire [1:0] v39; assign v39[1:0] = model_inp[79:78]; // 0.0
    wire [1:0] v40; assign v40[1:0] = model_inp[81:80]; // 0.0
    wire [1:0] v41; assign v41[1:0] = model_inp[83:82]; // 0.0
    wire [1:0] v42; assign v42[1:0] = model_inp[85:84]; // 0.0
    wire [1:0] v43; assign v43[1:0] = model_inp[87:86]; // 0.0
    wire [1:0] v44; assign v44[1:0] = model_inp[89:88]; // 0.0
    wire [1:0] v45; assign v45[1:0] = model_inp[91:90]; // 0.0
    wire [1:0] v46; assign v46[1:0] = model_inp[93:92]; // 0.0
    wire [1:0] v47; assign v47[1:0] = model_inp[95:94]; // 0.0
    wire [1:0] v48; assign v48[1:0] = model_inp[97:96]; // 0.0
    wire [1:0] v49; assign v49[1:0] = model_inp[99:98]; // 0.0
    wire [1:0] v50; assign v50[1:0] = model_inp[101:100]; // 0.0
    wire [1:0] v51; assign v51[1:0] = model_inp[103:102]; // 0.0
    wire [1:0] v52; assign v52[1:0] = model_inp[105:104]; // 0.0
    wire [1:0] v53; assign v53[1:0] = model_inp[107:106]; // 0.0
    wire [1:0] v54; assign v54[1:0] = model_inp[109:108]; // 0.0
    wire [1:0] v55; assign v55[1:0] = model_inp[111:110]; // 0.0
    wire [1:0] v56; assign v56[1:0] = model_inp[113:112]; // 0.0
    wire [1:0] v57; assign v57[1:0] = model_inp[115:114]; // 0.0
    wire [1:0] v58; assign v58[1:0] = model_inp[117:116]; // 0.0
    wire [1:0] v59; assign v59[1:0] = model_inp[119:118]; // 0.0
    wire [1:0] v60; assign v60[1:0] = v21[1:0]; // 0.0
    wire [2:0] v61; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_61 (v60[1:0], 1'b1, v61[2:0]); // 0.0
    wire [0:0] v62; assign v62[0:0] = v61[1:1]; // 0.0
    wire [1:0] v63; assign v63[1:0] = v14[1:0]; // 0.0
    wire [2:0] v64; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_64 (v63[1:0], 1'b1, v64[2:0]); // 0.0
    wire [0:0] v65; assign v65[0:0] = v64[1:1]; // 0.0
    wire [1:0] v66; assign v66[1:0] = v18[1:0]; // 0.0
    wire [2:0] v67; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_67 (v66[1:0], 1'b1, v67[2:0]); // 0.0
    wire [0:0] v68; assign v68[0:0] = v67[1:1]; // 0.0
    wire [1:0] v69; assign v69[1:0] = v20[1:0]; // 0.0
    wire [2:0] v70; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_70 (v69[1:0], 1'b1, v70[2:0]); // 0.0
    wire [0:0] v71; assign v71[0:0] = v70[1:1]; // 0.0
    wire [1:0] v72; assign v72[1:0] = v7[1:0]; // 0.0
    wire [2:0] v73; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_73 (v72[1:0], 1'b1, v73[2:0]); // 0.0
    wire [0:0] v74; assign v74[0:0] = v73[1:1]; // 0.0
    wire [1:0] v75; assign v75[1:0] = v22[1:0]; // 0.0
    wire [2:0] v76; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_76 (v75[1:0], 1'b1, v76[2:0]); // 0.0
    wire [0:0] v77; assign v77[0:0] = v76[1:1]; // 0.0
    wire [1:0] v78; assign v78[1:0] = v6[1:0]; // 0.0
    wire [2:0] v79; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_79 (v78[1:0], 1'b1, v79[2:0]); // 0.0
    wire [0:0] v80; assign v80[0:0] = v79[1:1]; // 0.0
    wire [1:0] v81; assign v81[1:0] = v17[1:0]; // 0.0
    wire [2:0] v82; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_82 (v81[1:0], 1'b1, v82[2:0]); // 0.0
    wire [0:0] v83; assign v83[0:0] = v82[1:1]; // 0.0
    wire [1:0] v84; assign v84[1:0] = v10[1:0]; // 0.0
    wire [2:0] v85; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_85 (v84[1:0], 1'b1, v85[2:0]); // 0.0
    wire [0:0] v86; assign v86[0:0] = v85[1:1]; // 0.0
    wire [1:0] v87; assign v87[1:0] = v19[1:0]; // 0.0
    wire [2:0] v88; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_88 (v87[1:0], 1'b1, v88[2:0]); // 0.0
    wire [0:0] v89; assign v89[0:0] = v88[1:1]; // 0.0
    wire [1:0] v90; assign v90[1:0] = v11[1:0]; // 0.0
    wire [2:0] v91; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_91 (v90[1:0], 1'b1, v91[2:0]); // 0.0
    wire [0:0] v92; assign v92[0:0] = v91[1:1]; // 0.0
    wire [1:0] v93; assign v93[1:0] = v23[1:0]; // 0.0
    wire [2:0] v94; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_94 (v93[1:0], 1'b1, v94[2:0]); // 0.0
    wire [0:0] v95; assign v95[0:0] = v94[1:1]; // 0.0
    wire [1:0] v96; assign v96[1:0] = v13[1:0]; // 0.0
    wire [2:0] v97; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_97 (v96[1:0], 1'b1, v97[2:0]); // 0.0
    wire [0:0] v98; assign v98[0:0] = v97[1:1]; // 0.0
    wire [1:0] v99; assign v99[1:0] = v12[1:0]; // 0.0
    wire [2:0] v100; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_100 (v99[1:0], 1'b1, v100[2:0]); // 0.0
    wire [0:0] v101; assign v101[0:0] = v100[1:1]; // 0.0
    wire [1:0] v102; assign v102[1:0] = v15[1:0]; // 0.0
    wire [2:0] v103; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_103 (v102[1:0], 1'b1, v103[2:0]); // 0.0
    wire [0:0] v104; assign v104[0:0] = v103[1:1]; // 0.0
    wire [1:0] v105; assign v105[1:0] = v9[1:0]; // 0.0
    wire [2:0] v106; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_106 (v105[1:0], 1'b1, v106[2:0]); // 0.0
    wire [0:0] v107; assign v107[0:0] = v106[1:1]; // 0.0
    wire [1:0] v108; assign v108[1:0] = v8[1:0]; // 0.0
    wire [2:0] v109; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_109 (v108[1:0], 1'b1, v109[2:0]); // 0.0
    wire [0:0] v110; assign v110[0:0] = v109[1:1]; // 0.0
    wire [1:0] v111; assign v111[1:0] = v16[1:0]; // 0.0
    wire [2:0] v112; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_112 (v111[1:0], 1'b1, v112[2:0]); // 0.0
    wire [0:0] v113; assign v113[0:0] = v112[1:1]; // 0.0
    wire [1:0] v114; assign v114[1:0] = v4[1:0]; // 0.0
    wire [2:0] v115; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_115 (v114[1:0], 1'b1, v115[2:0]); // 0.0
    wire [0:0] v116; assign v116[0:0] = v115[1:1]; // 0.0
    wire [1:0] v117; assign v117[1:0] = v3[1:0]; // 0.0
    wire [2:0] v118; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_118 (v117[1:0], 1'b1, v118[2:0]); // 0.0
    wire [0:0] v119; assign v119[0:0] = v118[1:1]; // 0.0
    wire [1:0] v120; assign v120[1:0] = v2[1:0]; // 0.0
    wire [2:0] v121; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_121 (v120[1:0], 1'b1, v121[2:0]); // 0.0
    wire [0:0] v122; assign v122[0:0] = v121[1:1]; // 0.0
    wire [1:0] v123; assign v123[1:0] = v0[1:0]; // 0.0
    wire [2:0] v124; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_124 (v123[1:0], 1'b1, v124[2:0]); // 0.0
    wire [0:0] v125; assign v125[0:0] = v124[1:1]; // 0.0
    wire [1:0] v126; assign v126[1:0] = v5[1:0]; // 0.0
    wire [2:0] v127; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_127 (v126[1:0], 1'b1, v127[2:0]); // 0.0
    wire [0:0] v128; assign v128[0:0] = v127[1:1]; // 0.0
    wire [1:0] v129; assign v129[1:0] = v1[1:0]; // 0.0
    wire [2:0] v130; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_130 (v129[1:0], 1'b1, v130[2:0]); // 0.0
    wire [0:0] v131; assign v131[0:0] = v130[1:1]; // 0.0
    wire [1:0] v132; assign v132[1:0] = v26[1:0]; // 0.0
    wire [2:0] v133; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_133 (v132[1:0], 1'b1, v133[2:0]); // 0.0
    wire [0:0] v134; assign v134[0:0] = v133[1:1]; // 0.0
    wire [1:0] v135; assign v135[1:0] = v28[1:0]; // 0.0
    wire [2:0] v136; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_136 (v135[1:0], 1'b1, v136[2:0]); // 0.0
    wire [0:0] v137; assign v137[0:0] = v136[1:1]; // 0.0
    wire [1:0] v138; assign v138[1:0] = v25[1:0]; // 0.0
    wire [2:0] v139; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_139 (v138[1:0], 1'b1, v139[2:0]); // 0.0
    wire [0:0] v140; assign v140[0:0] = v139[1:1]; // 0.0
    wire [1:0] v141; assign v141[1:0] = v27[1:0]; // 0.0
    wire [2:0] v142; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_142 (v141[1:0], 1'b1, v142[2:0]); // 0.0
    wire [0:0] v143; assign v143[0:0] = v142[1:1]; // 0.0
    wire [1:0] v144; assign v144[1:0] = v24[1:0]; // 0.0
    wire [2:0] v145; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_145 (v144[1:0], 1'b1, v145[2:0]); // 0.0
    wire [0:0] v146; assign v146[0:0] = v145[1:1]; // 0.0
    wire [1:0] v147; assign v147[1:0] = v29[1:0]; // 0.0
    wire [2:0] v148; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_148 (v147[1:0], 1'b1, v148[2:0]); // 0.0
    wire [0:0] v149; assign v149[0:0] = v148[1:1]; // 0.0
    wire [1:0] v150; assign v150[1:0] = v32[1:0]; // 0.0
    wire [2:0] v151; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_151 (v150[1:0], 1'b1, v151[2:0]); // 0.0
    wire [0:0] v152; assign v152[0:0] = v151[1:1]; // 0.0
    wire [1:0] v153; assign v153[1:0] = v30[1:0]; // 0.0
    wire [2:0] v154; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_154 (v153[1:0], 1'b1, v154[2:0]); // 0.0
    wire [0:0] v155; assign v155[0:0] = v154[1:1]; // 0.0
    wire [1:0] v156; assign v156[1:0] = v35[1:0]; // 0.0
    wire [2:0] v157; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_157 (v156[1:0], 1'b1, v157[2:0]); // 0.0
    wire [0:0] v158; assign v158[0:0] = v157[1:1]; // 0.0
    wire [1:0] v159; assign v159[1:0] = v33[1:0]; // 0.0
    wire [2:0] v160; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_160 (v159[1:0], 1'b1, v160[2:0]); // 0.0
    wire [0:0] v161; assign v161[0:0] = v160[1:1]; // 0.0
    wire [1:0] v162; assign v162[1:0] = v31[1:0]; // 0.0
    wire [2:0] v163; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_163 (v162[1:0], 1'b1, v163[2:0]); // 0.0
    wire [0:0] v164; assign v164[0:0] = v163[1:1]; // 0.0
    wire [1:0] v165; assign v165[1:0] = v34[1:0]; // 0.0
    wire [2:0] v166; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_166 (v165[1:0], 1'b1, v166[2:0]); // 0.0
    wire [0:0] v167; assign v167[0:0] = v166[1:1]; // 0.0
    wire [1:0] v168; assign v168[1:0] = v38[1:0]; // 0.0
    wire [2:0] v169; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_169 (v168[1:0], 1'b1, v169[2:0]); // 0.0
    wire [0:0] v170; assign v170[0:0] = v169[1:1]; // 0.0
    wire [1:0] v171; assign v171[1:0] = v36[1:0]; // 0.0
    wire [2:0] v172; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_172 (v171[1:0], 1'b1, v172[2:0]); // 0.0
    wire [0:0] v173; assign v173[0:0] = v172[1:1]; // 0.0
    wire [1:0] v174; assign v174[1:0] = v41[1:0]; // 0.0
    wire [2:0] v175; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_175 (v174[1:0], 1'b1, v175[2:0]); // 0.0
    wire [0:0] v176; assign v176[0:0] = v175[1:1]; // 0.0
    wire [1:0] v177; assign v177[1:0] = v39[1:0]; // 0.0
    wire [2:0] v178; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_178 (v177[1:0], 1'b1, v178[2:0]); // 0.0
    wire [0:0] v179; assign v179[0:0] = v178[1:1]; // 0.0
    wire [1:0] v180; assign v180[1:0] = v37[1:0]; // 0.0
    wire [2:0] v181; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_181 (v180[1:0], 1'b1, v181[2:0]); // 0.0
    wire [0:0] v182; assign v182[0:0] = v181[1:1]; // 0.0
    wire [1:0] v183; assign v183[1:0] = v40[1:0]; // 0.0
    wire [2:0] v184; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_184 (v183[1:0], 1'b1, v184[2:0]); // 0.0
    wire [0:0] v185; assign v185[0:0] = v184[1:1]; // 0.0
    wire [1:0] v186; assign v186[1:0] = v44[1:0]; // 0.0
    wire [2:0] v187; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_187 (v186[1:0], 1'b1, v187[2:0]); // 0.0
    wire [0:0] v188; assign v188[0:0] = v187[1:1]; // 0.0
    wire [1:0] v189; assign v189[1:0] = v42[1:0]; // 0.0
    wire [2:0] v190; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_190 (v189[1:0], 1'b1, v190[2:0]); // 0.0
    wire [0:0] v191; assign v191[0:0] = v190[1:1]; // 0.0
    wire [1:0] v192; assign v192[1:0] = v47[1:0]; // 0.0
    wire [2:0] v193; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_193 (v192[1:0], 1'b1, v193[2:0]); // 0.0
    wire [0:0] v194; assign v194[0:0] = v193[1:1]; // 0.0
    wire [1:0] v195; assign v195[1:0] = v45[1:0]; // 0.0
    wire [2:0] v196; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_196 (v195[1:0], 1'b1, v196[2:0]); // 0.0
    wire [0:0] v197; assign v197[0:0] = v196[1:1]; // 0.0
    wire [1:0] v198; assign v198[1:0] = v43[1:0]; // 0.0
    wire [2:0] v199; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_199 (v198[1:0], 1'b1, v199[2:0]); // 0.0
    wire [0:0] v200; assign v200[0:0] = v199[1:1]; // 0.0
    wire [1:0] v201; assign v201[1:0] = v46[1:0]; // 0.0
    wire [2:0] v202; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_202 (v201[1:0], 1'b1, v202[2:0]); // 0.0
    wire [0:0] v203; assign v203[0:0] = v202[1:1]; // 0.0
    wire [1:0] v204; assign v204[1:0] = v50[1:0]; // 0.0
    wire [2:0] v205; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_205 (v204[1:0], 1'b1, v205[2:0]); // 0.0
    wire [0:0] v206; assign v206[0:0] = v205[1:1]; // 0.0
    wire [1:0] v207; assign v207[1:0] = v48[1:0]; // 0.0
    wire [2:0] v208; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_208 (v207[1:0], 1'b1, v208[2:0]); // 0.0
    wire [0:0] v209; assign v209[0:0] = v208[1:1]; // 0.0
    wire [1:0] v210; assign v210[1:0] = v53[1:0]; // 0.0
    wire [2:0] v211; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_211 (v210[1:0], 1'b1, v211[2:0]); // 0.0
    wire [0:0] v212; assign v212[0:0] = v211[1:1]; // 0.0
    wire [1:0] v213; assign v213[1:0] = v51[1:0]; // 0.0
    wire [2:0] v214; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_214 (v213[1:0], 1'b1, v214[2:0]); // 0.0
    wire [0:0] v215; assign v215[0:0] = v214[1:1]; // 0.0
    wire [1:0] v216; assign v216[1:0] = v49[1:0]; // 0.0
    wire [2:0] v217; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_217 (v216[1:0], 1'b1, v217[2:0]); // 0.0
    wire [0:0] v218; assign v218[0:0] = v217[1:1]; // 0.0
    wire [1:0] v219; assign v219[1:0] = v52[1:0]; // 0.0
    wire [2:0] v220; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_220 (v219[1:0], 1'b1, v220[2:0]); // 0.0
    wire [0:0] v221; assign v221[0:0] = v220[1:1]; // 0.0
    wire [1:0] v222; assign v222[1:0] = v56[1:0]; // 0.0
    wire [2:0] v223; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_223 (v222[1:0], 1'b1, v223[2:0]); // 0.0
    wire [0:0] v224; assign v224[0:0] = v223[1:1]; // 0.0
    wire [1:0] v225; assign v225[1:0] = v54[1:0]; // 0.0
    wire [2:0] v226; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_226 (v225[1:0], 1'b1, v226[2:0]); // 0.0
    wire [0:0] v227; assign v227[0:0] = v226[1:1]; // 0.0
    wire [1:0] v228; assign v228[1:0] = v59[1:0]; // 0.0
    wire [2:0] v229; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_229 (v228[1:0], 1'b1, v229[2:0]); // 0.0
    wire [0:0] v230; assign v230[0:0] = v229[1:1]; // 0.0
    wire [1:0] v231; assign v231[1:0] = v57[1:0]; // 0.0
    wire [2:0] v232; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_232 (v231[1:0], 1'b1, v232[2:0]); // 0.0
    wire [0:0] v233; assign v233[0:0] = v232[1:1]; // 0.0
    wire [1:0] v234; assign v234[1:0] = v55[1:0]; // 0.0
    wire [2:0] v235; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_235 (v234[1:0], 1'b1, v235[2:0]); // 0.0
    wire [0:0] v236; assign v236[0:0] = v235[1:1]; // 0.0
    wire [1:0] v237; assign v237[1:0] = v58[1:0]; // 0.0
    wire [2:0] v238; shift_adder #(2, 1, 0, 0, 3, 0, 0) op_238 (v237[1:0], 1'b1, v238[2:0]); // 0.0
    wire [0:0] v239; assign v239[0:0] = v238[1:1]; // 0.0
    wire [3:0] v240; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_240 (v62[0:0], v65[0:0], v240[3:0]); // 1.0
    wire [1:0] v241; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_241 (v68[0:0], v71[0:0], v241[1:0]); // 1.0
    wire [2:0] v242; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_242 (v74[0:0], v77[0:0], v242[2:0]); // 1.0
    wire [1:0] v243; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_243 (v80[0:0], v83[0:0], v243[1:0]); // 1.0
    wire [1:0] v244; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_244 (v86[0:0], v89[0:0], v244[1:0]); // 1.0
    wire [1:0] v245; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_245 (v101[0:0], v104[0:0], v245[1:0]); // 1.0
    wire [3:0] v246; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_246 (v98[0:0], v107[0:0], v246[3:0]); // 1.0
    wire [1:0] v247; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_247 (v110[0:0], v77[0:0], v247[1:0]); // 1.0
    wire [1:0] v248; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_248 (v86[0:0], v71[0:0], v248[1:0]); // 1.0
    wire [1:0] v249; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_249 (v65[0:0], v107[0:0], v249[1:0]); // 1.0
    wire [1:0] v250; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_250 (v80[0:0], v68[0:0], v250[1:0]); // 1.0
    wire [1:0] v251; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_251 (v116[0:0], v98[0:0], v251[1:0]); // 1.0
    wire [3:0] v252; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_252 (v74[0:0], v119[0:0], v252[3:0]); // 1.0
    wire [1:0] v253; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_253 (v122[0:0], v113[0:0], v253[1:0]); // 1.0
    wire [1:0] v254; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_254 (v116[0:0], v65[0:0], v254[1:0]); // 1.0
    wire [1:0] v255; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_255 (v110[0:0], v119[0:0], v255[1:0]); // 1.0
    wire [1:0] v256; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_256 (v125[0:0], v101[0:0], v256[1:0]); // 1.0
    wire [1:0] v257; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_257 (v80[0:0], v107[0:0], v257[1:0]); // 1.0
    wire [1:0] v258; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_258 (v116[0:0], v65[0:0], v258[1:0]); // 1.0
    wire [1:0] v259; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_259 (v122[0:0], v101[0:0], v259[1:0]); // 1.0
    wire [2:0] v260; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_260 (v92[0:0], v125[0:0], v260[2:0]); // 1.0
    wire [1:0] v261; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_261 (v107[0:0], v86[0:0], v261[1:0]); // 1.0
    wire [1:0] v262; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_262 (v110[0:0], v98[0:0], v262[1:0]); // 1.0
    wire [2:0] v263; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_263 (v122[0:0], v86[0:0], v263[2:0]); // 1.0
    wire [3:0] v264; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_264 (v80[0:0], v74[0:0], v264[3:0]); // 1.0
    wire [2:0] v265; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_265 (v110[0:0], v131[0:0], v265[2:0]); // 1.0
    wire [1:0] v266; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_266 (v125[0:0], v119[0:0], v266[1:0]); // 1.0
    wire [1:0] v267; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_267 (v125[0:0], v110[0:0], v267[1:0]); // 1.0
    wire [2:0] v268; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_268 (v131[0:0], v113[0:0], v268[2:0]); // 1.0
    wire [1:0] v269; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_269 (v86[0:0], v128[0:0], v269[1:0]); // 1.0
    wire [1:0] v270; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_270 (v122[0:0], v74[0:0], v270[1:0]); // 1.0
    wire [2:0] v271; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_271 (v128[0:0], v110[0:0], v271[2:0]); // 1.0
    wire [1:0] v272; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_272 (v119[0:0], v116[0:0], v272[1:0]); // 1.0
    wire [2:0] v273; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_273 (v92[0:0], v131[0:0], v273[2:0]); // 1.0
    wire [1:0] v274; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_274 (v101[0:0], v104[0:0], v274[1:0]); // 1.0
    wire [1:0] v275; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_275 (v110[0:0], v83[0:0], v275[1:0]); // 1.0
    wire [1:0] v276; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_276 (v74[0:0], v80[0:0], v276[1:0]); // 1.0
    wire [2:0] v277; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_277 (v128[0:0], v65[0:0], v277[2:0]); // 1.0
    wire [1:0] v278; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_278 (v98[0:0], v74[0:0], v278[1:0]); // 1.0
    wire [1:0] v279; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_279 (v86[0:0], v71[0:0], v279[1:0]); // 1.0
    wire [1:0] v280; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_280 (v110[0:0], v68[0:0], v280[1:0]); // 1.0
    wire [2:0] v281; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_281 (v83[0:0], v80[0:0], v281[2:0]); // 1.0
    wire [1:0] v282; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_282 (v104[0:0], v113[0:0], v282[1:0]); // 1.0
    wire [1:0] v283; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_283 (v65[0:0], v89[0:0], v283[1:0]); // 1.0
    wire [1:0] v284; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_284 (v86[0:0], v80[0:0], v284[1:0]); // 1.0
    wire [1:0] v285; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_285 (v128[0:0], v116[0:0], v285[1:0]); // 1.0
    wire [2:0] v286; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_286 (v92[0:0], v71[0:0], v286[2:0]); // 1.0
    wire [1:0] v287; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_287 (v89[0:0], v98[0:0], v287[1:0]); // 1.0
    wire [1:0] v288; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_288 (v80[0:0], v65[0:0], v288[1:0]); // 1.0
    wire [1:0] v289; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_289 (v113[0:0], v92[0:0], v289[1:0]); // 1.0
    wire [3:0] v290; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_290 (v74[0:0], v122[0:0], v290[3:0]); // 1.0
    wire [1:0] v291; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_291 (v107[0:0], v86[0:0], v291[1:0]); // 1.0
    wire [1:0] v292; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_292 (v128[0:0], v110[0:0], v292[1:0]); // 1.0
    wire [1:0] v293; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_293 (v116[0:0], v110[0:0], v293[1:0]); // 1.0
    wire [1:0] v294; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_294 (v80[0:0], v107[0:0], v294[1:0]); // 1.0
    wire [1:0] v295; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_295 (v92[0:0], v128[0:0], v295[1:0]); // 1.0
    wire [1:0] v296; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_296 (v80[0:0], v122[0:0], v296[1:0]); // 1.0
    wire [2:0] v297; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_297 (v92[0:0], v125[0:0], v297[2:0]); // 1.0
    wire [2:0] v298; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_298 (v83[0:0], v74[0:0], v298[2:0]); // 1.0
    wire [1:0] v299; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_299 (v68[0:0], v62[0:0], v299[1:0]); // 1.0
    wire [1:0] v300; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_300 (v65[0:0], v95[0:0], v300[1:0]); // 1.0
    wire [1:0] v301; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_301 (v98[0:0], v101[0:0], v301[1:0]); // 1.0
    wire [1:0] v302; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_302 (v77[0:0], v107[0:0], v302[1:0]); // 1.0
    wire [1:0] v303; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_303 (v62[0:0], v77[0:0], v303[1:0]); // 1.0
    wire [2:0] v304; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_304 (v83[0:0], v134[0:0], v304[2:0]); // 1.0
    wire [2:0] v305; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_305 (v98[0:0], v137[0:0], v305[2:0]); // 1.0
    wire [1:0] v306; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_306 (v140[0:0], v89[0:0], v306[1:0]); // 1.0
    wire [1:0] v307; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_307 (v71[0:0], v140[0:0], v307[1:0]); // 1.0
    wire [1:0] v308; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_308 (v65[0:0], v146[0:0], v308[1:0]); // 1.0
    wire [1:0] v309; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_309 (v113[0:0], v119[0:0], v309[1:0]); // 1.0
    wire [2:0] v310; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_310 (v95[0:0], v98[0:0], v310[2:0]); // 1.0
    wire [1:0] v311; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_311 (v101[0:0], v146[0:0], v311[1:0]); // 1.0
    wire [1:0] v312; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_312 (v113[0:0], v134[0:0], v312[1:0]); // 1.0
    wire [1:0] v313; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_313 (v146[0:0], v143[0:0], v313[1:0]); // 1.0
    wire [1:0] v314; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_314 (v65[0:0], v137[0:0], v314[1:0]); // 1.0
    wire [1:0] v315; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_315 (v71[0:0], v149[0:0], v315[1:0]); // 1.0
    wire [1:0] v316; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_316 (v89[0:0], v68[0:0], v316[1:0]); // 1.0
    wire [1:0] v317; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_317 (v68[0:0], v62[0:0], v317[1:0]); // 1.0
    wire [2:0] v318; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_318 (v95[0:0], v101[0:0], v318[2:0]); // 1.0
    wire [1:0] v319; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_319 (v101[0:0], v71[0:0], v319[1:0]); // 1.0
    wire [1:0] v320; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_320 (v113[0:0], v134[0:0], v320[1:0]); // 1.0
    wire [1:0] v321; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_321 (v77[0:0], v83[0:0], v321[1:0]); // 1.0
    wire [1:0] v322; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_322 (v137[0:0], v104[0:0], v322[1:0]); // 1.0
    wire [3:0] v323; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_323 (v104[0:0], v110[0:0], v323[3:0]); // 1.0
    wire [1:0] v324; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_324 (v101[0:0], v65[0:0], v324[1:0]); // 1.0
    wire [1:0] v325; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_325 (v125[0:0], v92[0:0], v325[1:0]); // 1.0
    wire [3:0] v326; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_326 (v143[0:0], v71[0:0], v326[3:0]); // 1.0
    wire [1:0] v327; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_327 (v146[0:0], v134[0:0], v327[1:0]); // 1.0
    wire [1:0] v328; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_328 (v101[0:0], v95[0:0], v328[1:0]); // 1.0
    wire [1:0] v329; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_329 (v113[0:0], v140[0:0], v329[1:0]); // 1.0
    wire [1:0] v330; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_330 (v77[0:0], v152[0:0], v330[1:0]); // 1.0
    wire [1:0] v331; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_331 (v71[0:0], v155[0:0], v331[1:0]); // 1.0
    wire [1:0] v332; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_332 (v146[0:0], v143[0:0], v332[1:0]); // 1.0
    wire [2:0] v333; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_333 (v149[0:0], v68[0:0], v333[2:0]); // 1.0
    wire [1:0] v334; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_334 (v143[0:0], v137[0:0], v334[1:0]); // 1.0
    wire [1:0] v335; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_335 (v134[0:0], v164[0:0], v335[1:0]); // 1.0
    wire [1:0] v336; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_336 (v167[0:0], v62[0:0], v336[1:0]); // 1.0
    wire [1:0] v337; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_337 (v68[0:0], v155[0:0], v337[1:0]); // 1.0
    wire [2:0] v338; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_338 (v95[0:0], v152[0:0], v338[2:0]); // 1.0
    wire [1:0] v339; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_339 (v68[0:0], v134[0:0], v339[1:0]); // 1.0
    wire [2:0] v340; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_340 (v89[0:0], v167[0:0], v340[2:0]); // 1.0
    wire [1:0] v341; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_341 (v77[0:0], v152[0:0], v341[1:0]); // 1.0
    wire [1:0] v342; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_342 (v137[0:0], v95[0:0], v342[1:0]); // 1.0
    wire [3:0] v343; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_343 (v89[0:0], v104[0:0], v343[3:0]); // 1.0
    wire [1:0] v344; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_344 (v71[0:0], v104[0:0], v344[1:0]); // 1.0
    wire [3:0] v345; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_345 (v161[0:0], v134[0:0], v345[3:0]); // 1.0
    wire [1:0] v346; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_346 (v155[0:0], v152[0:0], v346[1:0]); // 1.0
    wire [1:0] v347; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_347 (v68[0:0], v149[0:0], v347[1:0]); // 1.0
    wire [1:0] v348; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_348 (v77[0:0], v164[0:0], v348[1:0]); // 1.0
    wire [3:0] v349; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_349 (v140[0:0], v62[0:0], v349[3:0]); // 1.0
    wire [1:0] v350; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_350 (v71[0:0], v167[0:0], v350[1:0]); // 1.0
    wire [1:0] v351; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_351 (v134[0:0], v62[0:0], v351[1:0]); // 1.0
    wire [1:0] v352; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_352 (v164[0:0], v140[0:0], v352[1:0]); // 1.0
    wire [2:0] v353; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_353 (v149[0:0], v89[0:0], v353[2:0]); // 1.0
    wire [1:0] v354; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_354 (v155[0:0], v161[0:0], v354[1:0]); // 1.0
    wire [1:0] v355; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_355 (v134[0:0], v158[0:0], v355[1:0]); // 1.0
    wire [1:0] v356; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_356 (v140[0:0], v146[0:0], v356[1:0]); // 1.0
    wire [3:0] v357; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_357 (v110[0:0], v128[0:0], v357[3:0]); // 1.0
    wire [1:0] v358; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_358 (v137[0:0], v170[0:0], v358[1:0]); // 1.0
    wire [1:0] v359; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_359 (v134[0:0], v173[0:0], v359[1:0]); // 1.0
    wire [1:0] v360; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_360 (v155[0:0], v161[0:0], v360[1:0]); // 1.0
    wire [2:0] v361; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_361 (v158[0:0], v146[0:0], v361[2:0]); // 1.0
    wire [1:0] v362; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_362 (v161[0:0], v167[0:0], v362[1:0]); // 1.0
    wire [1:0] v363; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_363 (v152[0:0], v182[0:0], v363[1:0]); // 1.0
    wire [3:0] v364; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_364 (v179[0:0], v152[0:0], v364[3:0]); // 1.0
    wire [1:0] v365; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_365 (v173[0:0], v170[0:0], v365[1:0]); // 1.0
    wire [2:0] v366; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_366 (v140[0:0], v185[0:0], v366[2:0]); // 1.0
    wire [1:0] v367; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_367 (v146[0:0], v158[0:0], v367[1:0]); // 1.0
    wire [1:0] v368; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_368 (v137[0:0], v182[0:0], v368[1:0]); // 1.0
    wire [1:0] v369; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_369 (v146[0:0], v152[0:0], v369[1:0]); // 1.0
    wire [1:0] v370; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_370 (v137[0:0], v170[0:0], v370[1:0]); // 1.0
    wire [1:0] v371; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_371 (v167[0:0], v149[0:0], v371[1:0]); // 1.0
    wire [2:0] v372; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_372 (v149[0:0], v170[0:0], v372[2:0]); // 1.0
    wire [1:0] v373; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_373 (v182[0:0], v164[0:0], v373[1:0]); // 1.0
    wire [3:0] v374; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_374 (v164[0:0], v143[0:0], v374[3:0]); // 1.0
    wire [1:0] v375; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_375 (v134[0:0], v185[0:0], v375[1:0]); // 1.0
    wire [1:0] v376; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_376 (v152[0:0], v143[0:0], v376[1:0]); // 1.0
    wire [1:0] v377; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_377 (v146[0:0], v173[0:0], v377[1:0]); // 1.0
    wire [2:0] v378; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_378 (v158[0:0], v140[0:0], v378[2:0]); // 1.0
    wire [1:0] v379; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_379 (v173[0:0], v179[0:0], v379[1:0]); // 1.0
    wire [1:0] v380; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_380 (v152[0:0], v176[0:0], v380[1:0]); // 1.0
    wire [1:0] v381; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_381 (v164[0:0], v155[0:0], v381[1:0]); // 1.0
    wire [1:0] v382; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_382 (v167[0:0], v188[0:0], v382[1:0]); // 1.0
    wire [1:0] v383; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_383 (v152[0:0], v191[0:0], v383[1:0]); // 1.0
    wire [1:0] v384; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_384 (v173[0:0], v179[0:0], v384[1:0]); // 1.0
    wire [2:0] v385; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_385 (v176[0:0], v155[0:0], v385[2:0]); // 1.0
    wire [1:0] v386; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_386 (v179[0:0], v185[0:0], v386[1:0]); // 1.0
    wire [1:0] v387; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_387 (v170[0:0], v200[0:0], v387[1:0]); // 1.0
    wire [3:0] v388; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_388 (v197[0:0], v170[0:0], v388[3:0]); // 1.0
    wire [1:0] v389; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_389 (v191[0:0], v188[0:0], v389[1:0]); // 1.0
    wire [2:0] v390; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_390 (v164[0:0], v203[0:0], v390[2:0]); // 1.0
    wire [1:0] v391; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_391 (v155[0:0], v176[0:0], v391[1:0]); // 1.0
    wire [1:0] v392; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_392 (v167[0:0], v200[0:0], v392[1:0]); // 1.0
    wire [3:0] v393; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_393 (v182[0:0], v161[0:0], v393[3:0]); // 1.0
    wire [1:0] v394; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_394 (v152[0:0], v203[0:0], v394[1:0]); // 1.0
    wire [1:0] v395; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_395 (v167[0:0], v188[0:0], v395[1:0]); // 1.0
    wire [1:0] v396; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_396 (v170[0:0], v161[0:0], v396[1:0]); // 1.0
    wire [1:0] v397; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_397 (v155[0:0], v191[0:0], v397[1:0]); // 1.0
    wire [1:0] v398; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_398 (v155[0:0], v170[0:0], v398[1:0]); // 1.0
    wire [1:0] v399; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_399 (v185[0:0], v158[0:0], v399[1:0]); // 1.0
    wire [2:0] v400; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_400 (v158[0:0], v188[0:0], v400[2:0]); // 1.0
    wire [1:0] v401; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_401 (v200[0:0], v182[0:0], v401[1:0]); // 1.0
    wire [2:0] v402; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_402 (v176[0:0], v164[0:0], v402[2:0]); // 1.0
    wire [1:0] v403; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_403 (v191[0:0], v197[0:0], v403[1:0]); // 1.0
    wire [1:0] v404; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_404 (v170[0:0], v194[0:0], v404[1:0]); // 1.0
    wire [1:0] v405; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_405 (v182[0:0], v173[0:0], v405[1:0]); // 1.0
    wire [1:0] v406; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_406 (v203[0:0], v161[0:0], v406[1:0]); // 1.0
    wire [1:0] v407; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_407 (v185[0:0], v143[0:0], v407[1:0]); // 1.0
    wire [1:0] v408; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_408 (v185[0:0], v206[0:0], v408[1:0]); // 1.0
    wire [1:0] v409; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_409 (v170[0:0], v209[0:0], v409[1:0]); // 1.0
    wire [1:0] v410; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_410 (v191[0:0], v197[0:0], v410[1:0]); // 1.0
    wire [2:0] v411; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_411 (v194[0:0], v173[0:0], v411[2:0]); // 1.0
    wire [1:0] v412; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_412 (v197[0:0], v203[0:0], v412[1:0]); // 1.0
    wire [1:0] v413; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_413 (v188[0:0], v218[0:0], v413[1:0]); // 1.0
    wire [3:0] v414; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_414 (v215[0:0], v188[0:0], v414[3:0]); // 1.0
    wire [1:0] v415; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_415 (v209[0:0], v206[0:0], v415[1:0]); // 1.0
    wire [2:0] v416; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_416 (v182[0:0], v221[0:0], v416[2:0]); // 1.0
    wire [1:0] v417; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_417 (v173[0:0], v194[0:0], v417[1:0]); // 1.0
    wire [1:0] v418; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_418 (v185[0:0], v218[0:0], v418[1:0]); // 1.0
    wire [3:0] v419; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_419 (v200[0:0], v179[0:0], v419[3:0]); // 1.0
    wire [1:0] v420; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_420 (v170[0:0], v221[0:0], v420[1:0]); // 1.0
    wire [1:0] v421; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_421 (v185[0:0], v206[0:0], v421[1:0]); // 1.0
    wire [1:0] v422; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_422 (v188[0:0], v179[0:0], v422[1:0]); // 1.0
    wire [1:0] v423; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_423 (v173[0:0], v209[0:0], v423[1:0]); // 1.0
    wire [1:0] v424; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_424 (v173[0:0], v188[0:0], v424[1:0]); // 1.0
    wire [1:0] v425; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_425 (v203[0:0], v176[0:0], v425[1:0]); // 1.0
    wire [2:0] v426; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_426 (v176[0:0], v206[0:0], v426[2:0]); // 1.0
    wire [1:0] v427; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_427 (v218[0:0], v200[0:0], v427[1:0]); // 1.0
    wire [2:0] v428; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_428 (v194[0:0], v182[0:0], v428[2:0]); // 1.0
    wire [1:0] v429; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_429 (v209[0:0], v215[0:0], v429[1:0]); // 1.0
    wire [1:0] v430; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_430 (v188[0:0], v212[0:0], v430[1:0]); // 1.0
    wire [1:0] v431; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_431 (v200[0:0], v191[0:0], v431[1:0]); // 1.0
    wire [1:0] v432; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_432 (v221[0:0], v179[0:0], v432[1:0]); // 1.0
    wire [1:0] v433; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_433 (v203[0:0], v224[0:0], v433[1:0]); // 1.0
    wire [1:0] v434; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_434 (v188[0:0], v227[0:0], v434[1:0]); // 1.0
    wire [1:0] v435; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_435 (v209[0:0], v215[0:0], v435[1:0]); // 1.0
    wire [2:0] v436; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_436 (v212[0:0], v191[0:0], v436[2:0]); // 1.0
    wire [1:0] v437; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_437 (v215[0:0], v221[0:0], v437[1:0]); // 1.0
    wire [1:0] v438; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_438 (v206[0:0], v236[0:0], v438[1:0]); // 1.0
    wire [1:0] v439; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_439 (v203[0:0], v236[0:0], v439[1:0]); // 1.0
    wire [3:0] v440; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_440 (v218[0:0], v197[0:0], v440[3:0]); // 1.0
    wire [1:0] v441; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_441 (v188[0:0], v239[0:0], v441[1:0]); // 1.0
    wire [1:0] v442; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_442 (v203[0:0], v224[0:0], v442[1:0]); // 1.0
    wire [1:0] v443; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_443 (v206[0:0], v197[0:0], v443[1:0]); // 1.0
    wire [1:0] v444; shift_adder #(1, 1, 0, 0, 2, 1, 1) op_444 (v191[0:0], v227[0:0], v444[1:0]); // 1.0
    wire [3:0] v445; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_445 (v233[0:0], v206[0:0], v445[3:0]); // 1.0
    wire [1:0] v446; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_446 (v227[0:0], v224[0:0], v446[1:0]); // 1.0
    wire [2:0] v447; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_447 (v200[0:0], v239[0:0], v447[2:0]); // 1.0
    wire [1:0] v448; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_448 (v191[0:0], v212[0:0], v448[1:0]); // 1.0
    wire [1:0] v449; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_449 (v191[0:0], v206[0:0], v449[1:0]); // 1.0
    wire [1:0] v450; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_450 (v221[0:0], v194[0:0], v450[1:0]); // 1.0
    wire [2:0] v451; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_451 (v194[0:0], v224[0:0], v451[2:0]); // 1.0
    wire [1:0] v452; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_452 (v236[0:0], v218[0:0], v452[1:0]); // 1.0
    wire [1:0] v453; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_453 (v239[0:0], v197[0:0], v453[1:0]); // 1.0
    wire [2:0] v454; shift_adder #(1, 1, 0, 0, 3, 2, 0) op_454 (v212[0:0], v200[0:0], v454[2:0]); // 1.0
    wire [1:0] v455; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_455 (v227[0:0], v233[0:0], v455[1:0]); // 1.0
    wire [1:0] v456; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_456 (v206[0:0], v230[0:0], v456[1:0]); // 1.0
    wire [1:0] v457; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_457 (v218[0:0], v209[0:0], v457[1:0]); // 1.0
    wire [1:0] v458; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_458 (v209[0:0], v221[0:0], v458[1:0]); // 1.0
    wire [2:0] v459; shift_adder #(1, 1, 0, 0, 3, -1, 1) op_459 (v218[0:0], v230[0:0], v459[2:0]); // 1.0
    wire [1:0] v460; shift_adder #(1, 1, 0, 0, 2, 1, 0) op_460 (v224[0:0], v206[0:0], v460[1:0]); // 1.0
    wire [1:0] v461; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_461 (v227[0:0], v236[0:0], v461[1:0]); // 1.0
    wire [1:0] v462; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_462 (v233[0:0], v239[0:0], v462[1:0]); // 1.0
    wire [1:0] v463; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_463 (v212[0:0], v236[0:0], v463[1:0]); // 1.0
    wire [1:0] v464; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_464 (v206[0:0], v224[0:0], v464[1:0]); // 1.0
    wire [1:0] v465; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_465 (v230[0:0], v215[0:0], v465[1:0]); // 1.0
    wire [2:0] v466; shift_adder #(1, 1, 0, 0, 3, 2, 1) op_466 (v221[0:0], v239[0:0], v466[2:0]); // 1.0
    wire [3:0] v467; shift_adder #(1, 1, 0, 0, 4, -2, 1) op_467 (v215[0:0], v215[0:0], v467[3:0]); // 1.0
    wire [1:0] v468; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_468 (v209[0:0], v221[0:0], v468[1:0]); // 1.0
    wire [2:0] v469; shift_adder #(1, 1, 0, 0, 3, -2, 0) op_469 (v218[0:0], v230[0:0], v469[2:0]); // 1.0
    wire [1:0] v470; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_470 (v227[0:0], v212[0:0], v470[1:0]); // 1.0
    wire [1:0] v471; shift_adder #(1, 1, 0, 0, 2, 0, 1) op_471 (v233[0:0], v209[0:0], v471[1:0]); // 1.0
    wire [1:0] v472; shift_adder #(1, 1, 0, 0, 2, -1, 0) op_472 (v224[0:0], v239[0:0], v472[1:0]); // 1.0
    wire [1:0] v473; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_473 (v206[0:0], v224[0:0], v473[1:0]); // 1.0
    wire [4:0] v474; shift_adder #(4, 2, 1, 0, 5, 1, 0) op_474 (v240[3:0], v241[1:0], v474[4:0]); // 2.0
    wire [3:0] v475; shift_adder #(2, 2, 0, 1, 4, 0, 0) op_475 (v243[1:0], v244[1:0], v475[3:0]); // 2.0
    wire [2:0] v476; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_476 (v98[0:0], v245[1:0], v476[2:0]); // 2.0
    wire [4:0] v477; shift_adder #(2, 4, 1, 1, 5, 1, 0) op_477 (v244[1:0], v246[3:0], v477[4:0]); // 2.0
    wire [3:0] v478; shift_adder #(2, 2, 0, 0, 4, 1, 0) op_478 (v248[1:0], v249[1:0], v478[3:0]); // 2.0
    wire [2:0] v479; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_479 (v113[0:0], v250[1:0], v479[2:0]); // 2.0
    wire [4:0] v480; shift_adder #(2, 4, 1, 1, 5, 1, 0) op_480 (v251[1:0], v252[3:0], v480[4:0]); // 2.0
    wire [3:0] v481; shift_adder #(2, 2, 0, 0, 4, 1, 0) op_481 (v254[1:0], v255[1:0], v481[3:0]); // 2.0
    wire [2:0] v482; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_482 (v86[0:0], v256[1:0], v482[2:0]); // 2.0
    wire [2:0] v483; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_483 (v74[0:0], v257[1:0], v483[2:0]); // 2.0
    wire [1:0] v484; shift_adder #(2, 1, 1, 0, 2, 0, 1) op_484 (v258[1:0], v128[0:0], v484[1:0]); // 2.0
    wire [4:0] v485; shift_adder #(3, 2, 1, 0, 5, 1, 0) op_485 (v260[2:0], v261[1:0], v485[4:0]); // 2.0
    wire [2:0] v486; shift_adder #(1, 2, 0, 1, 3, -1, 1) op_486 (v119[0:0], v262[1:0], v486[2:0]); // 2.0
    wire [2:0] v487; shift_adder #(3, 1, 1, 0, 3, 1, 1) op_487 (v263[2:0], v116[0:0], v487[2:0]); // 2.0
    wire [4:0] v488; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_488 (v264[3:0], v265[2:0], v488[4:0]); // 2.0
    wire [2:0] v489; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_489 (v131[0:0], v266[1:0], v489[2:0]); // 2.0
    wire [2:0] v490; shift_adder #(2, 1, 0, 0, 3, 0, 1) op_490 (v267[1:0], v83[0:0], v490[2:0]); // 2.0
    wire [2:0] v491; shift_adder #(1, 2, 0, 1, 3, 1, 1) op_491 (v104[0:0], v259[1:0], v491[2:0]); // 2.0
    wire [2:0] v492; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_492 (v92[0:0], v268[2:0], v492[2:0]); // 2.0
    wire [2:0] v493; shift_adder #(2, 2, 0, 0, 3, 1, 0) op_493 (v254[1:0], v269[1:0], v493[2:0]); // 2.0
    wire [2:0] v494; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_494 (v107[0:0], v270[1:0], v494[2:0]); // 2.0
    wire [4:0] v495; shift_adder #(3, 2, 1, 0, 5, 1, 0) op_495 (v271[2:0], v272[1:0], v495[4:0]); // 2.0
    wire [4:0] v496; shift_adder #(3, 2, 0, 1, 5, 2, 0) op_496 (v273[2:0], v256[1:0], v496[4:0]); // 2.0
    wire [2:0] v497; shift_adder #(2, 2, 1, 0, 3, 0, 0) op_497 (v258[1:0], v274[1:0], v497[2:0]); // 2.0
    wire [2:0] v498; shift_adder #(2, 2, 0, 0, 3, 0, 0) op_498 (v261[1:0], v253[1:0], v498[2:0]); // 2.0
    wire [3:0] v499; shift_adder #(2, 2, 0, 0, 4, -1, 1) op_499 (v275[1:0], v276[1:0], v499[3:0]); // 2.0
    wire [3:0] v500; shift_adder #(2, 3, 0, 0, 4, 0, 0) op_500 (v261[1:0], v277[2:0], v500[3:0]); // 2.0
    wire [3:0] v501; shift_adder #(2, 1, 0, 0, 4, 3, 1) op_501 (v278[1:0], v74[0:0], v501[3:0]); // 2.0
    wire [1:0] v502; shift_adder #(2, 1, 1, 0, 2, 0, 1) op_502 (v279[1:0], v92[0:0], v502[1:0]); // 2.0
    wire [4:0] v503; shift_adder #(3, 2, 1, 0, 5, 1, 0) op_503 (v281[2:0], v282[1:0], v503[4:0]); // 2.0
    wire [2:0] v504; shift_adder #(1, 2, 0, 1, 3, -1, 1) op_504 (v107[0:0], v283[1:0], v504[2:0]); // 2.0
    wire [2:0] v505; shift_adder #(2, 1, 0, 0, 3, 2, 1) op_505 (v284[1:0], v110[0:0], v505[2:0]); // 2.0
    wire [3:0] v506; shift_adder #(2, 2, 1, 0, 4, 0, 0) op_506 (v266[1:0], v285[1:0], v506[3:0]); // 2.0
    wire [3:0] v507; shift_adder #(2, 3, 0, 0, 4, 0, 0) op_507 (v282[1:0], v286[2:0], v507[3:0]); // 2.0
    wire [2:0] v508; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_508 (v83[0:0], v242[2:0], v508[2:0]); // 2.0
    wire [3:0] v509; shift_adder #(2, 1, 0, 0, 4, 3, 1) op_509 (v287[1:0], v98[0:0], v509[3:0]); // 2.0
    wire [2:0] v510; shift_adder #(1, 2, 0, 1, 3, 1, 1) op_510 (v62[0:0], v280[1:0], v510[2:0]); // 2.0
    wire [2:0] v511; shift_adder #(2, 1, 0, 0, 3, 0, 1) op_511 (v288[1:0], v95[0:0], v511[2:0]); // 2.0
    wire [2:0] v512; shift_adder #(2, 2, 0, 0, 3, 1, 0) op_512 (v248[1:0], v289[1:0], v512[2:0]); // 2.0
    wire [4:0] v513; shift_adder #(4, 2, 1, 0, 5, 2, 0) op_513 (v290[3:0], v291[1:0], v513[4:0]); // 2.0
    wire [3:0] v514; shift_adder #(3, 2, 1, 0, 4, -1, 1) op_514 (v263[2:0], v293[1:0], v514[3:0]); // 2.0
    wire [3:0] v515; shift_adder #(2, 2, 0, 0, 4, -1, 0) op_515 (v294[1:0], v295[1:0], v515[3:0]); // 2.0
    wire [4:0] v516; shift_adder #(2, 1, 1, 0, 5, 3, 1) op_516 (v292[1:0], v80[0:0], v516[4:0]); // 2.0
    wire [3:0] v517; shift_adder #(3, 2, 1, 0, 4, 0, 0) op_517 (v297[2:0], v272[1:0], v517[3:0]); // 2.0
    wire [1:0] v518; shift_adder #(1, 2, 0, 0, 2, 0, 1) op_518 (v131[0:0], v291[1:0], v518[1:0]); // 2.0
    wire [4:0] v519; shift_adder #(3, 2, 0, 1, 5, 2, 0) op_519 (v298[2:0], v250[1:0], v519[4:0]); // 2.0
    wire [2:0] v520; shift_adder #(2, 2, 1, 0, 3, 0, 0) op_520 (v279[1:0], v299[1:0], v520[2:0]); // 2.0
    wire [2:0] v521; shift_adder #(2, 2, 0, 0, 3, 0, 0) op_521 (v282[1:0], v247[1:0], v521[2:0]); // 2.0
    wire [3:0] v522; shift_adder #(2, 2, 0, 0, 4, -1, 1) op_522 (v300[1:0], v301[1:0], v522[3:0]); // 2.0
    wire [2:0] v523; shift_adder #(2, 1, 1, 0, 3, 1, 1) op_523 (v302[1:0], v83[0:0], v523[2:0]); // 2.0
    wire [3:0] v524; shift_adder #(3, 2, 0, 1, 4, 0, 0) op_524 (v286[2:0], v245[1:0], v524[3:0]); // 2.0
    wire [3:0] v525; shift_adder #(2, 3, 0, 0, 4, 0, 0) op_525 (v303[1:0], v304[2:0], v525[3:0]); // 2.0
    wire [2:0] v526; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_526 (v95[0:0], v305[2:0], v526[2:0]); // 2.0
    wire [3:0] v527; shift_adder #(2, 1, 0, 0, 4, 3, 1) op_527 (v306[1:0], v89[0:0], v527[3:0]); // 2.0
    wire [2:0] v528; shift_adder #(1, 2, 0, 1, 3, 1, 1) op_528 (v143[0:0], v308[1:0], v528[2:0]); // 2.0
    wire [2:0] v529; shift_adder #(2, 1, 1, 0, 3, 1, 1) op_529 (v309[1:0], v92[0:0], v529[2:0]); // 2.0
    wire [3:0] v530; shift_adder #(3, 2, 0, 1, 4, 0, 0) op_530 (v277[2:0], v257[1:0], v530[3:0]); // 2.0
    wire [4:0] v531; shift_adder #(3, 2, 0, 1, 5, 2, 0) op_531 (v310[2:0], v311[1:0], v531[4:0]); // 2.0
    wire [2:0] v532; shift_adder #(2, 2, 1, 0, 3, 0, 0) op_532 (v312[1:0], v313[1:0], v532[2:0]); // 2.0
    wire [2:0] v533; shift_adder #(2, 2, 0, 0, 3, 0, 0) op_533 (v303[1:0], v314[1:0], v533[2:0]); // 2.0
    wire [3:0] v534; shift_adder #(2, 2, 0, 0, 4, -1, 1) op_534 (v315[1:0], v316[1:0], v534[3:0]); // 2.0
    wire [1:0] v535; shift_adder #(2, 1, 1, 0, 2, 0, 1) op_535 (v312[1:0], v83[0:0], v535[1:0]); // 2.0
    wire [2:0] v536; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_536 (v89[0:0], v317[1:0], v536[2:0]); // 2.0
    wire [4:0] v537; shift_adder #(3, 2, 1, 0, 5, 1, 0) op_537 (v318[2:0], v303[1:0], v537[4:0]); // 2.0
    wire [2:0] v538; shift_adder #(1, 2, 0, 1, 3, -1, 1) op_538 (v104[0:0], v307[1:0], v538[2:0]); // 2.0
    wire [2:0] v539; shift_adder #(2, 1, 0, 0, 3, 0, 1) op_539 (v319[1:0], v149[0:0], v539[2:0]); // 2.0
    wire [2:0] v540; shift_adder #(2, 2, 0, 0, 3, 1, 0) op_540 (v320[1:0], v321[1:0], v540[2:0]); // 2.0
    wire [2:0] v541; shift_adder #(2, 1, 1, 0, 3, 1, 1) op_541 (v322[1:0], v95[0:0], v541[2:0]); // 2.0
    wire [2:0] v542; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_542 (v77[0:0], v311[1:0], v542[2:0]); // 2.0
    wire [3:0] v543; shift_adder #(3, 2, 0, 1, 4, 0, 0) op_543 (v304[2:0], v317[1:0], v543[3:0]); // 2.0
    wire [4:0] v544; shift_adder #(4, 2, 1, 0, 5, 1, 0) op_544 (v323[3:0], v324[1:0], v544[4:0]); // 2.0
    wire [3:0] v545; shift_adder #(2, 2, 0, 1, 4, 0, 0) op_545 (v325[1:0], v251[1:0], v545[3:0]); // 2.0
    wire [4:0] v546; shift_adder #(4, 2, 1, 0, 5, 1, 0) op_546 (v326[3:0], v327[1:0], v546[4:0]); // 2.0
    wire [3:0] v547; shift_adder #(2, 2, 0, 1, 4, 0, 0) op_547 (v328[1:0], v329[1:0], v547[3:0]); // 2.0
    wire [1:0] v548; shift_adder #(2, 1, 1, 0, 2, 0, 1) op_548 (v330[1:0], v95[0:0], v548[1:0]); // 2.0
    wire [2:0] v549; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_549 (v140[0:0], v332[1:0], v549[2:0]); // 2.0
    wire [4:0] v550; shift_adder #(3, 2, 1, 0, 5, 1, 0) op_550 (v333[2:0], v334[1:0], v550[4:0]); // 2.0
    wire [2:0] v551; shift_adder #(1, 2, 0, 1, 3, -1, 1) op_551 (v62[0:0], v335[1:0], v551[2:0]); // 2.0
    wire [2:0] v552; shift_adder #(2, 1, 1, 0, 3, 1, 1) op_552 (v336[1:0], v149[0:0], v552[2:0]); // 2.0
    wire [2:0] v553; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_553 (v137[0:0], v337[1:0], v553[2:0]); // 2.0
    wire [3:0] v554; shift_adder #(3, 2, 0, 1, 4, 0, 0) op_554 (v338[2:0], v332[1:0], v554[3:0]); // 2.0
    wire [2:0] v555; shift_adder #(2, 1, 0, 0, 3, 0, 1) op_555 (v339[1:0], v158[0:0], v555[2:0]); // 2.0
    wire [2:0] v556; shift_adder #(1, 2, 0, 1, 3, 1, 1) op_556 (v161[0:0], v331[1:0], v556[2:0]); // 2.0
    wire [2:0] v557; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_557 (v149[0:0], v340[2:0], v557[2:0]); // 2.0
    wire [2:0] v558; shift_adder #(2, 2, 0, 0, 3, 1, 0) op_558 (v341[1:0], v342[1:0], v558[2:0]); // 2.0
    wire [4:0] v559; shift_adder #(2, 4, 1, 1, 5, 1, 0) op_559 (v329[1:0], v343[3:0], v559[4:0]); // 2.0
    wire [3:0] v560; shift_adder #(2, 2, 0, 0, 4, 1, 0) op_560 (v320[1:0], v344[1:0], v560[3:0]); // 2.0
    wire [4:0] v561; shift_adder #(4, 2, 1, 0, 5, 1, 0) op_561 (v345[3:0], v346[1:0], v561[4:0]); // 2.0
    wire [3:0] v562; shift_adder #(2, 2, 0, 1, 4, 0, 0) op_562 (v347[1:0], v348[1:0], v562[3:0]); // 2.0
    wire [4:0] v563; shift_adder #(2, 4, 1, 1, 5, 1, 0) op_563 (v348[1:0], v349[3:0], v563[4:0]); // 2.0
    wire [3:0] v564; shift_adder #(2, 2, 0, 0, 4, 1, 0) op_564 (v341[1:0], v351[1:0], v564[3:0]); // 2.0
    wire [3:0] v565; shift_adder #(2, 3, 0, 0, 4, 0, 0) op_565 (v334[1:0], v338[2:0], v565[3:0]); // 2.0
    wire [3:0] v566; shift_adder #(2, 1, 0, 0, 4, 3, 1) op_566 (v352[1:0], v140[0:0], v566[3:0]); // 2.0
    wire [4:0] v567; shift_adder #(3, 2, 0, 1, 5, 2, 0) op_567 (v353[2:0], v337[1:0], v567[4:0]); // 2.0
    wire [2:0] v568; shift_adder #(2, 2, 1, 0, 3, 0, 0) op_568 (v330[1:0], v354[1:0], v568[2:0]); // 2.0
    wire [2:0] v569; shift_adder #(2, 2, 0, 0, 3, 0, 0) op_569 (v334[1:0], v350[1:0], v569[2:0]); // 2.0
    wire [3:0] v570; shift_adder #(2, 2, 0, 0, 4, -1, 1) op_570 (v355[1:0], v356[1:0], v570[3:0]); // 2.0
    wire [3:0] v571; shift_adder #(4, 1, 1, 0, 4, 2, 1) op_571 (v357[3:0], v131[0:0], v571[3:0]); // 2.0
    wire [3:0] v572; shift_adder #(2, 4, 0, 1, 4, -1, 1) op_572 (v272[1:0], v264[3:0], v572[3:0]); // 2.0
    wire [1:0] v573; shift_adder #(2, 1, 1, 0, 2, 0, 1) op_573 (v358[1:0], v149[0:0], v573[1:0]); // 2.0
    wire [2:0] v574; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_574 (v164[0:0], v360[1:0], v574[2:0]); // 2.0
    wire [4:0] v575; shift_adder #(3, 2, 1, 0, 5, 1, 0) op_575 (v361[2:0], v362[1:0], v575[4:0]); // 2.0
    wire [2:0] v576; shift_adder #(1, 2, 0, 1, 3, -1, 1) op_576 (v143[0:0], v363[1:0], v576[2:0]); // 2.0
    wire [4:0] v577; shift_adder #(4, 2, 1, 0, 5, 1, 0) op_577 (v364[3:0], v365[1:0], v577[4:0]); // 2.0
    wire [3:0] v578; shift_adder #(2, 2, 0, 1, 4, 0, 0) op_578 (v367[1:0], v368[1:0], v578[3:0]); // 2.0
    wire [2:0] v579; shift_adder #(2, 1, 0, 0, 3, 0, 1) op_579 (v369[1:0], v176[0:0], v579[2:0]); // 2.0
    wire [2:0] v580; shift_adder #(1, 2, 0, 1, 3, 1, 1) op_580 (v179[0:0], v359[1:0], v580[2:0]); // 2.0
    wire [2:0] v581; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_581 (v158[0:0], v366[2:0], v581[2:0]); // 2.0
    wire [2:0] v582; shift_adder #(2, 2, 0, 0, 3, 1, 0) op_582 (v370[1:0], v371[1:0], v582[2:0]); // 2.0
    wire [3:0] v583; shift_adder #(2, 3, 0, 0, 4, 0, 0) op_583 (v362[1:0], v372[2:0], v583[3:0]); // 2.0
    wire [3:0] v584; shift_adder #(2, 1, 0, 0, 4, 3, 1) op_584 (v373[1:0], v164[0:0], v584[3:0]); // 2.0
    wire [4:0] v585; shift_adder #(2, 4, 1, 1, 5, 1, 0) op_585 (v368[1:0], v374[3:0], v585[4:0]); // 2.0
    wire [3:0] v586; shift_adder #(2, 2, 0, 0, 4, 1, 0) op_586 (v370[1:0], v376[1:0], v586[3:0]); // 2.0
    wire [2:0] v587; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_587 (v167[0:0], v377[1:0], v587[2:0]); // 2.0
    wire [4:0] v588; shift_adder #(3, 2, 0, 1, 5, 2, 0) op_588 (v378[2:0], v377[1:0], v588[4:0]); // 2.0
    wire [2:0] v589; shift_adder #(2, 2, 1, 0, 3, 0, 0) op_589 (v358[1:0], v379[1:0], v589[2:0]); // 2.0
    wire [2:0] v590; shift_adder #(2, 2, 0, 0, 3, 0, 0) op_590 (v362[1:0], v375[1:0], v590[2:0]); // 2.0
    wire [3:0] v591; shift_adder #(2, 2, 0, 0, 4, -1, 1) op_591 (v380[1:0], v381[1:0], v591[3:0]); // 2.0
    wire [1:0] v592; shift_adder #(2, 1, 1, 0, 2, 0, 1) op_592 (v382[1:0], v158[0:0], v592[1:0]); // 2.0
    wire [2:0] v593; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_593 (v182[0:0], v384[1:0], v593[2:0]); // 2.0
    wire [4:0] v594; shift_adder #(3, 2, 1, 0, 5, 1, 0) op_594 (v385[2:0], v386[1:0], v594[4:0]); // 2.0
    wire [2:0] v595; shift_adder #(1, 2, 0, 1, 3, -1, 1) op_595 (v161[0:0], v387[1:0], v595[2:0]); // 2.0
    wire [4:0] v596; shift_adder #(4, 2, 1, 0, 5, 1, 0) op_596 (v388[3:0], v389[1:0], v596[4:0]); // 2.0
    wire [3:0] v597; shift_adder #(2, 2, 0, 1, 4, 0, 0) op_597 (v391[1:0], v392[1:0], v597[3:0]); // 2.0
    wire [4:0] v598; shift_adder #(2, 4, 1, 1, 5, 1, 0) op_598 (v392[1:0], v393[3:0], v598[4:0]); // 2.0
    wire [3:0] v599; shift_adder #(2, 2, 0, 0, 4, 1, 0) op_599 (v395[1:0], v396[1:0], v599[3:0]); // 2.0
    wire [2:0] v600; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_600 (v185[0:0], v397[1:0], v600[2:0]); // 2.0
    wire [2:0] v601; shift_adder #(2, 1, 0, 0, 3, 0, 1) op_601 (v398[1:0], v194[0:0], v601[2:0]); // 2.0
    wire [2:0] v602; shift_adder #(1, 2, 0, 1, 3, 1, 1) op_602 (v197[0:0], v383[1:0], v602[2:0]); // 2.0
    wire [2:0] v603; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_603 (v176[0:0], v390[2:0], v603[2:0]); // 2.0
    wire [2:0] v604; shift_adder #(2, 2, 0, 0, 3, 1, 0) op_604 (v395[1:0], v399[1:0], v604[2:0]); // 2.0
    wire [3:0] v605; shift_adder #(2, 3, 0, 0, 4, 0, 0) op_605 (v386[1:0], v400[2:0], v605[3:0]); // 2.0
    wire [3:0] v606; shift_adder #(2, 1, 0, 0, 4, 3, 1) op_606 (v401[1:0], v182[0:0], v606[3:0]); // 2.0
    wire [4:0] v607; shift_adder #(3, 2, 0, 1, 5, 2, 0) op_607 (v402[2:0], v397[1:0], v607[4:0]); // 2.0
    wire [2:0] v608; shift_adder #(2, 2, 1, 0, 3, 0, 0) op_608 (v382[1:0], v403[1:0], v608[2:0]); // 2.0
    wire [2:0] v609; shift_adder #(2, 2, 0, 0, 3, 0, 0) op_609 (v386[1:0], v394[1:0], v609[2:0]); // 2.0
    wire [3:0] v610; shift_adder #(2, 2, 0, 0, 4, -1, 1) op_610 (v404[1:0], v405[1:0], v610[3:0]); // 2.0
    wire [2:0] v611; shift_adder #(2, 1, 1, 0, 3, 1, 1) op_611 (v406[1:0], v176[0:0], v611[2:0]); // 2.0
    wire [3:0] v612; shift_adder #(3, 2, 0, 1, 4, 0, 0) op_612 (v400[2:0], v384[1:0], v612[3:0]); // 2.0
    wire [2:0] v613; shift_adder #(2, 1, 1, 0, 3, 1, 1) op_613 (v407[1:0], v158[0:0], v613[2:0]); // 2.0
    wire [3:0] v614; shift_adder #(3, 2, 0, 1, 4, 0, 0) op_614 (v372[2:0], v360[1:0], v614[3:0]); // 2.0
    wire [1:0] v615; shift_adder #(2, 1, 1, 0, 2, 0, 1) op_615 (v408[1:0], v176[0:0], v615[1:0]); // 2.0
    wire [2:0] v616; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_616 (v200[0:0], v410[1:0], v616[2:0]); // 2.0
    wire [4:0] v617; shift_adder #(3, 2, 1, 0, 5, 1, 0) op_617 (v411[2:0], v412[1:0], v617[4:0]); // 2.0
    wire [2:0] v618; shift_adder #(1, 2, 0, 1, 3, -1, 1) op_618 (v179[0:0], v413[1:0], v618[2:0]); // 2.0
    wire [4:0] v619; shift_adder #(4, 2, 1, 0, 5, 1, 0) op_619 (v414[3:0], v415[1:0], v619[4:0]); // 2.0
    wire [3:0] v620; shift_adder #(2, 2, 0, 1, 4, 0, 0) op_620 (v417[1:0], v418[1:0], v620[3:0]); // 2.0
    wire [4:0] v621; shift_adder #(2, 4, 1, 1, 5, 1, 0) op_621 (v418[1:0], v419[3:0], v621[4:0]); // 2.0
    wire [3:0] v622; shift_adder #(2, 2, 0, 0, 4, 1, 0) op_622 (v421[1:0], v422[1:0], v622[3:0]); // 2.0
    wire [2:0] v623; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_623 (v203[0:0], v423[1:0], v623[2:0]); // 2.0
    wire [2:0] v624; shift_adder #(2, 1, 0, 0, 3, 0, 1) op_624 (v424[1:0], v212[0:0], v624[2:0]); // 2.0
    wire [2:0] v625; shift_adder #(1, 2, 0, 1, 3, 1, 1) op_625 (v215[0:0], v409[1:0], v625[2:0]); // 2.0
    wire [2:0] v626; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_626 (v194[0:0], v416[2:0], v626[2:0]); // 2.0
    wire [2:0] v627; shift_adder #(2, 2, 0, 0, 3, 1, 0) op_627 (v421[1:0], v425[1:0], v627[2:0]); // 2.0
    wire [3:0] v628; shift_adder #(2, 3, 0, 0, 4, 0, 0) op_628 (v412[1:0], v426[2:0], v628[3:0]); // 2.0
    wire [3:0] v629; shift_adder #(2, 1, 0, 0, 4, 3, 1) op_629 (v427[1:0], v200[0:0], v629[3:0]); // 2.0
    wire [4:0] v630; shift_adder #(3, 2, 0, 1, 5, 2, 0) op_630 (v428[2:0], v423[1:0], v630[4:0]); // 2.0
    wire [2:0] v631; shift_adder #(2, 2, 1, 0, 3, 0, 0) op_631 (v408[1:0], v429[1:0], v631[2:0]); // 2.0
    wire [2:0] v632; shift_adder #(2, 2, 0, 0, 3, 0, 0) op_632 (v412[1:0], v420[1:0], v632[2:0]); // 2.0
    wire [3:0] v633; shift_adder #(2, 2, 0, 0, 4, -1, 1) op_633 (v430[1:0], v431[1:0], v633[3:0]); // 2.0
    wire [2:0] v634; shift_adder #(2, 1, 1, 0, 3, 1, 1) op_634 (v432[1:0], v194[0:0], v634[2:0]); // 2.0
    wire [3:0] v635; shift_adder #(3, 2, 0, 1, 4, 0, 0) op_635 (v426[2:0], v410[1:0], v635[3:0]); // 2.0
    wire [1:0] v636; shift_adder #(2, 1, 1, 0, 2, 0, 1) op_636 (v433[1:0], v194[0:0], v636[1:0]); // 2.0
    wire [2:0] v637; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_637 (v218[0:0], v435[1:0], v637[2:0]); // 2.0
    wire [4:0] v638; shift_adder #(3, 2, 1, 0, 5, 1, 0) op_638 (v436[2:0], v437[1:0], v638[4:0]); // 2.0
    wire [2:0] v639; shift_adder #(1, 2, 0, 1, 3, -1, 1) op_639 (v197[0:0], v438[1:0], v639[2:0]); // 2.0
    wire [4:0] v640; shift_adder #(2, 4, 1, 1, 5, 1, 0) op_640 (v439[1:0], v440[3:0], v640[4:0]); // 2.0
    wire [3:0] v641; shift_adder #(2, 2, 0, 0, 4, 1, 0) op_641 (v442[1:0], v443[1:0], v641[3:0]); // 2.0
    wire [2:0] v642; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_642 (v221[0:0], v444[1:0], v642[2:0]); // 2.0
    wire [4:0] v643; shift_adder #(4, 2, 1, 0, 5, 1, 0) op_643 (v445[3:0], v446[1:0], v643[4:0]); // 2.0
    wire [3:0] v644; shift_adder #(2, 2, 0, 1, 4, 0, 0) op_644 (v448[1:0], v439[1:0], v644[3:0]); // 2.0
    wire [2:0] v645; shift_adder #(2, 1, 0, 0, 3, 0, 1) op_645 (v449[1:0], v230[0:0], v645[2:0]); // 2.0
    wire [2:0] v646; shift_adder #(1, 2, 0, 1, 3, 1, 1) op_646 (v233[0:0], v434[1:0], v646[2:0]); // 2.0
    wire [2:0] v647; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_647 (v212[0:0], v447[2:0], v647[2:0]); // 2.0
    wire [2:0] v648; shift_adder #(2, 2, 0, 0, 3, 1, 0) op_648 (v442[1:0], v450[1:0], v648[2:0]); // 2.0
    wire [3:0] v649; shift_adder #(2, 3, 0, 0, 4, 0, 0) op_649 (v437[1:0], v451[2:0], v649[3:0]); // 2.0
    wire [3:0] v650; shift_adder #(2, 1, 0, 0, 4, 3, 1) op_650 (v452[1:0], v218[0:0], v650[3:0]); // 2.0
    wire [2:0] v651; shift_adder #(2, 1, 1, 0, 3, 1, 1) op_651 (v453[1:0], v212[0:0], v651[2:0]); // 2.0
    wire [3:0] v652; shift_adder #(3, 2, 0, 1, 4, 0, 0) op_652 (v451[2:0], v435[1:0], v652[3:0]); // 2.0
    wire [4:0] v653; shift_adder #(3, 2, 0, 1, 5, 2, 0) op_653 (v454[2:0], v444[1:0], v653[4:0]); // 2.0
    wire [2:0] v654; shift_adder #(2, 2, 1, 0, 3, 0, 0) op_654 (v433[1:0], v455[1:0], v654[2:0]); // 2.0
    wire [2:0] v655; shift_adder #(2, 2, 0, 0, 3, 0, 0) op_655 (v437[1:0], v441[1:0], v655[2:0]); // 2.0
    wire [3:0] v656; shift_adder #(2, 2, 0, 0, 4, -1, 1) op_656 (v456[1:0], v457[1:0], v656[3:0]); // 2.0
    wire [1:0] v657; shift_adder #(2, 1, 1, 0, 2, 0, 1) op_657 (v458[1:0], v239[0:0], v657[1:0]); // 2.0
    wire [4:0] v658; shift_adder #(3, 2, 1, 0, 5, 1, 0) op_658 (v459[2:0], v460[1:0], v658[4:0]); // 2.0
    wire [1:0] v659; shift_adder #(1, 2, 0, 0, 2, 0, 1) op_659 (v233[0:0], v461[1:0], v659[1:0]); // 2.0
    wire [3:0] v660; shift_adder #(3, 2, 1, 0, 4, 0, 0) op_660 (v459[2:0], v463[1:0], v660[3:0]); // 2.0
    wire [2:0] v661; shift_adder #(1, 2, 0, 1, 3, -1, 1) op_661 (v236[0:0], v464[1:0], v661[2:0]); // 2.0
    wire [3:0] v662; shift_adder #(2, 2, 1, 0, 4, 0, 0) op_662 (v465[1:0], v462[1:0], v662[3:0]); // 2.0
    wire [2:0] v663; shift_adder #(2, 2, 1, 1, 3, 0, 0) op_663 (v458[1:0], v464[1:0], v663[2:0]); // 2.0
    wire [4:0] v664; shift_adder #(3, 4, 1, 1, 5, 1, 0) op_664 (v466[2:0], v467[3:0], v664[4:0]); // 2.0
    wire [2:0] v665; shift_adder #(2, 1, 0, 0, 3, -1, 0) op_665 (v468[1:0], v224[0:0], v665[2:0]); // 2.0
    wire [3:0] v666; shift_adder #(4, 2, 1, 0, 4, 0, 1) op_666 (v467[3:0], v470[1:0], v666[3:0]); // 2.0
    wire [2:0] v667; shift_adder #(2, 1, 1, 0, 3, 1, 1) op_667 (v471[1:0], v230[0:0], v667[2:0]); // 2.0
    wire [2:0] v668; shift_adder #(2, 2, 0, 0, 3, 1, 0) op_668 (v468[1:0], v473[1:0], v668[2:0]); // 2.0
    wire [3:0] v669; shift_adder #(3, 2, 0, 0, 4, 1, 0) op_669 (v469[2:0], v462[1:0], v669[3:0]); // 2.0
    wire [4:0] v670; shift_adder #(5, 3, 1, 1, 5, 2, 1) op_670 (v474[4:0], v242[2:0], v670[4:0]); // 3.0
    wire [2:0] v671; shift_adder #(1, 3, 0, 1, 3, 0, 0) op_671 (v95[0:0], v476[2:0], v671[2:0]); // 3.0
    wire [4:0] v672; shift_adder #(5, 2, 1, 0, 5, 1, 1) op_672 (v477[4:0], v247[1:0], v672[4:0]); // 3.0
    wire [4:0] v673; shift_adder #(4, 3, 0, 1, 5, 1, 1) op_673 (v478[3:0], v479[2:0], v673[4:0]); // 3.0
    wire [4:0] v674; shift_adder #(5, 2, 1, 0, 5, 1, 1) op_674 (v480[4:0], v253[1:0], v674[4:0]); // 3.0
    wire [4:0] v675; shift_adder #(4, 3, 0, 1, 5, 1, 1) op_675 (v481[3:0], v482[2:0], v675[4:0]); // 3.0
    wire [2:0] v676; shift_adder #(1, 3, 0, 1, 3, 0, 0) op_676 (v83[0:0], v483[2:0], v676[2:0]); // 3.0
    wire [2:0] v677; shift_adder #(2, 2, 1, 1, 3, 0, 1) op_677 (v484[1:0], v259[1:0], v677[2:0]); // 3.0
    wire [2:0] v678; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_678 (v104[0:0], v486[2:0], v678[2:0]); // 3.0
    wire [4:0] v679; shift_adder #(3, 5, 1, 1, 5, 0, 0) op_679 (v487[2:0], v488[4:0], v679[4:0]); // 3.0
    wire [2:0] v680; shift_adder #(1, 3, 0, 1, 3, 0, 0) op_680 (v92[0:0], v489[2:0], v680[2:0]); // 3.0
    wire [3:0] v681; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_681 (v483[2:0], v490[2:0], v681[3:0]); // 3.0
    wire [4:0] v682; shift_adder #(3, 3, 1, 0, 5, -1, 0) op_682 (v492[2:0], v493[2:0], v682[4:0]); // 3.0
    wire [4:0] v683; shift_adder #(3, 5, 1, 1, 5, 0, 0) op_683 (v494[2:0], v495[4:0], v683[4:0]); // 3.0
    wire [4:0] v684; shift_adder #(5, 3, 1, 1, 5, 1, 0) op_684 (v496[4:0], v497[2:0], v684[4:0]); // 3.0
    wire [4:0] v685; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_685 (v498[2:0], v499[3:0], v685[4:0]); // 3.0
    wire [4:0] v686; shift_adder #(4, 3, 0, 1, 5, 0, 1) op_686 (v500[3:0], v492[2:0], v686[4:0]); // 3.0
    wire [4:0] v687; shift_adder #(4, 2, 1, 1, 5, 2, 1) op_687 (v501[3:0], v262[1:0], v687[4:0]); // 3.0
    wire [2:0] v688; shift_adder #(2, 2, 1, 1, 3, 0, 1) op_688 (v502[1:0], v280[1:0], v688[2:0]); // 3.0
    wire [2:0] v689; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_689 (v62[0:0], v504[2:0], v689[2:0]); // 3.0
    wire [3:0] v690; shift_adder #(3, 3, 1, 1, 4, 1, 1) op_690 (v505[2:0], v494[2:0], v690[3:0]); // 3.0
    wire [4:0] v691; shift_adder #(4, 3, 0, 1, 5, 0, 1) op_691 (v507[3:0], v508[2:0], v691[4:0]); // 3.0
    wire [4:0] v692; shift_adder #(4, 2, 1, 1, 5, 2, 1) op_692 (v509[3:0], v283[1:0], v692[4:0]); // 3.0
    wire [3:0] v693; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_693 (v476[2:0], v511[2:0], v693[3:0]); // 3.0
    wire [4:0] v694; shift_adder #(3, 3, 1, 0, 5, -1, 0) op_694 (v508[2:0], v512[2:0], v694[4:0]); // 3.0
    wire [5:0] v695; shift_adder #(5, 2, 1, 1, 6, 1, 1) op_695 (v513[4:0], v292[1:0], v695[5:0]); // 3.0
    wire [4:0] v696; shift_adder #(3, 4, 1, 1, 5, -1, 0) op_696 (v489[2:0], v514[3:0], v696[4:0]); // 3.0
    wire [4:0] v697; shift_adder #(2, 5, 0, 1, 5, -1, 0) op_697 (v296[1:0], v516[4:0], v697[4:0]); // 3.0
    wire [3:0] v698; shift_adder #(4, 2, 1, 1, 4, 0, 1) op_698 (v517[3:0], v518[1:0], v698[3:0]); // 3.0
    wire [4:0] v699; shift_adder #(5, 3, 1, 1, 5, 1, 0) op_699 (v519[4:0], v520[2:0], v699[4:0]); // 3.0
    wire [4:0] v700; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_700 (v521[2:0], v522[3:0], v700[4:0]); // 3.0
    wire [3:0] v701; shift_adder #(3, 3, 1, 1, 4, 0, 1) op_701 (v523[2:0], v479[2:0], v701[3:0]); // 3.0
    wire [4:0] v702; shift_adder #(4, 3, 0, 1, 5, 0, 1) op_702 (v525[3:0], v526[2:0], v702[4:0]); // 3.0
    wire [4:0] v703; shift_adder #(4, 2, 1, 1, 5, 2, 1) op_703 (v527[3:0], v307[1:0], v703[4:0]); // 3.0
    wire [3:0] v704; shift_adder #(3, 3, 1, 1, 4, 0, 1) op_704 (v529[2:0], v482[2:0], v704[3:0]); // 3.0
    wire [4:0] v705; shift_adder #(5, 3, 1, 1, 5, 1, 0) op_705 (v531[4:0], v532[2:0], v705[4:0]); // 3.0
    wire [4:0] v706; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_706 (v533[2:0], v534[3:0], v706[4:0]); // 3.0
    wire [2:0] v707; shift_adder #(2, 2, 1, 1, 3, 0, 1) op_707 (v535[1:0], v308[1:0], v707[2:0]); // 3.0
    wire [2:0] v708; shift_adder #(1, 3, 0, 1, 3, 0, 0) op_708 (v149[0:0], v536[2:0], v708[2:0]); // 3.0
    wire [2:0] v709; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_709 (v143[0:0], v538[2:0], v709[2:0]); // 3.0
    wire [3:0] v710; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_710 (v536[2:0], v539[2:0], v710[3:0]); // 3.0
    wire [4:0] v711; shift_adder #(3, 3, 1, 0, 5, -1, 0) op_711 (v526[2:0], v540[2:0], v711[4:0]); // 3.0
    wire [3:0] v712; shift_adder #(3, 3, 1, 1, 4, 0, 1) op_712 (v541[2:0], v542[2:0], v712[3:0]); // 3.0
    wire [4:0] v713; shift_adder #(5, 3, 1, 1, 5, 2, 1) op_713 (v544[4:0], v268[2:0], v713[4:0]); // 3.0
    wire [4:0] v714; shift_adder #(5, 3, 1, 1, 5, 2, 1) op_714 (v546[4:0], v305[2:0], v714[4:0]); // 3.0
    wire [2:0] v715; shift_adder #(2, 2, 1, 1, 3, 0, 1) op_715 (v548[1:0], v331[1:0], v715[2:0]); // 3.0
    wire [2:0] v716; shift_adder #(1, 3, 0, 1, 3, 0, 0) op_716 (v158[0:0], v549[2:0], v716[2:0]); // 3.0
    wire [2:0] v717; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_717 (v161[0:0], v551[2:0], v717[2:0]); // 3.0
    wire [3:0] v718; shift_adder #(3, 3, 1, 1, 4, 0, 1) op_718 (v552[2:0], v553[2:0], v718[3:0]); // 3.0
    wire [3:0] v719; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_719 (v549[2:0], v555[2:0], v719[3:0]); // 3.0
    wire [4:0] v720; shift_adder #(3, 3, 1, 0, 5, -1, 0) op_720 (v557[2:0], v558[2:0], v720[4:0]); // 3.0
    wire [4:0] v721; shift_adder #(5, 2, 1, 0, 5, 1, 1) op_721 (v559[4:0], v314[1:0], v721[4:0]); // 3.0
    wire [4:0] v722; shift_adder #(4, 3, 0, 1, 5, 1, 1) op_722 (v560[3:0], v542[2:0], v722[4:0]); // 3.0
    wire [4:0] v723; shift_adder #(5, 3, 1, 1, 5, 2, 1) op_723 (v561[4:0], v340[2:0], v723[4:0]); // 3.0
    wire [4:0] v724; shift_adder #(5, 2, 1, 0, 5, 1, 1) op_724 (v563[4:0], v350[1:0], v724[4:0]); // 3.0
    wire [4:0] v725; shift_adder #(4, 3, 0, 1, 5, 1, 1) op_725 (v564[3:0], v553[2:0], v725[4:0]); // 3.0
    wire [4:0] v726; shift_adder #(4, 3, 0, 1, 5, 0, 1) op_726 (v565[3:0], v557[2:0], v726[4:0]); // 3.0
    wire [4:0] v727; shift_adder #(4, 2, 1, 1, 5, 2, 1) op_727 (v566[3:0], v335[1:0], v727[4:0]); // 3.0
    wire [4:0] v728; shift_adder #(5, 3, 1, 1, 5, 1, 0) op_728 (v567[4:0], v568[2:0], v728[4:0]); // 3.0
    wire [4:0] v729; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_729 (v569[2:0], v570[3:0], v729[4:0]); // 3.0
    wire [2:0] v730; shift_adder #(2, 2, 1, 1, 3, 1, 1) op_730 (v518[1:0], v270[1:0], v730[2:0]); // 3.0
    wire [4:0] v731; shift_adder #(4, 4, 1, 1, 5, -1, 0) op_731 (v571[3:0], v572[3:0], v731[4:0]); // 3.0
    wire [2:0] v732; shift_adder #(2, 2, 1, 1, 3, 0, 1) op_732 (v573[1:0], v359[1:0], v732[2:0]); // 3.0
    wire [2:0] v733; shift_adder #(1, 3, 0, 1, 3, 0, 0) op_733 (v176[0:0], v574[2:0], v733[2:0]); // 3.0
    wire [2:0] v734; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_734 (v179[0:0], v576[2:0], v734[2:0]); // 3.0
    wire [4:0] v735; shift_adder #(5, 3, 1, 1, 5, 2, 1) op_735 (v577[4:0], v366[2:0], v735[4:0]); // 3.0
    wire [3:0] v736; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_736 (v574[2:0], v579[2:0], v736[3:0]); // 3.0
    wire [4:0] v737; shift_adder #(3, 3, 1, 0, 5, -1, 0) op_737 (v581[2:0], v582[2:0], v737[4:0]); // 3.0
    wire [4:0] v738; shift_adder #(4, 3, 0, 1, 5, 0, 1) op_738 (v583[3:0], v581[2:0], v738[4:0]); // 3.0
    wire [4:0] v739; shift_adder #(4, 2, 1, 1, 5, 2, 1) op_739 (v584[3:0], v363[1:0], v739[4:0]); // 3.0
    wire [4:0] v740; shift_adder #(5, 2, 1, 0, 5, 1, 1) op_740 (v585[4:0], v375[1:0], v740[4:0]); // 3.0
    wire [4:0] v741; shift_adder #(4, 3, 0, 1, 5, 1, 1) op_741 (v586[3:0], v587[2:0], v741[4:0]); // 3.0
    wire [4:0] v742; shift_adder #(5, 3, 1, 1, 5, 1, 0) op_742 (v588[4:0], v589[2:0], v742[4:0]); // 3.0
    wire [4:0] v743; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_743 (v590[2:0], v591[3:0], v743[4:0]); // 3.0
    wire [2:0] v744; shift_adder #(2, 2, 1, 1, 3, 0, 1) op_744 (v592[1:0], v383[1:0], v744[2:0]); // 3.0
    wire [2:0] v745; shift_adder #(1, 3, 0, 1, 3, 0, 0) op_745 (v194[0:0], v593[2:0], v745[2:0]); // 3.0
    wire [2:0] v746; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_746 (v197[0:0], v595[2:0], v746[2:0]); // 3.0
    wire [4:0] v747; shift_adder #(5, 3, 1, 1, 5, 2, 1) op_747 (v596[4:0], v390[2:0], v747[4:0]); // 3.0
    wire [4:0] v748; shift_adder #(5, 2, 1, 0, 5, 1, 1) op_748 (v598[4:0], v394[1:0], v748[4:0]); // 3.0
    wire [4:0] v749; shift_adder #(4, 3, 0, 1, 5, 1, 1) op_749 (v599[3:0], v600[2:0], v749[4:0]); // 3.0
    wire [3:0] v750; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_750 (v593[2:0], v601[2:0], v750[3:0]); // 3.0
    wire [4:0] v751; shift_adder #(3, 3, 1, 0, 5, -1, 0) op_751 (v603[2:0], v604[2:0], v751[4:0]); // 3.0
    wire [4:0] v752; shift_adder #(4, 3, 0, 1, 5, 0, 1) op_752 (v605[3:0], v603[2:0], v752[4:0]); // 3.0
    wire [4:0] v753; shift_adder #(4, 2, 1, 1, 5, 2, 1) op_753 (v606[3:0], v387[1:0], v753[4:0]); // 3.0
    wire [4:0] v754; shift_adder #(5, 3, 1, 1, 5, 1, 0) op_754 (v607[4:0], v608[2:0], v754[4:0]); // 3.0
    wire [4:0] v755; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_755 (v609[2:0], v610[3:0], v755[4:0]); // 3.0
    wire [3:0] v756; shift_adder #(3, 3, 1, 1, 4, 0, 1) op_756 (v611[2:0], v600[2:0], v756[3:0]); // 3.0
    wire [3:0] v757; shift_adder #(3, 3, 1, 1, 4, 0, 1) op_757 (v613[2:0], v587[2:0], v757[3:0]); // 3.0
    wire [2:0] v758; shift_adder #(2, 2, 1, 1, 3, 0, 1) op_758 (v615[1:0], v409[1:0], v758[2:0]); // 3.0
    wire [2:0] v759; shift_adder #(1, 3, 0, 1, 3, 0, 0) op_759 (v212[0:0], v616[2:0], v759[2:0]); // 3.0
    wire [2:0] v760; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_760 (v215[0:0], v618[2:0], v760[2:0]); // 3.0
    wire [4:0] v761; shift_adder #(5, 3, 1, 1, 5, 2, 1) op_761 (v619[4:0], v416[2:0], v761[4:0]); // 3.0
    wire [4:0] v762; shift_adder #(5, 2, 1, 0, 5, 1, 1) op_762 (v621[4:0], v420[1:0], v762[4:0]); // 3.0
    wire [4:0] v763; shift_adder #(4, 3, 0, 1, 5, 1, 1) op_763 (v622[3:0], v623[2:0], v763[4:0]); // 3.0
    wire [3:0] v764; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_764 (v616[2:0], v624[2:0], v764[3:0]); // 3.0
    wire [4:0] v765; shift_adder #(3, 3, 1, 0, 5, -1, 0) op_765 (v626[2:0], v627[2:0], v765[4:0]); // 3.0
    wire [4:0] v766; shift_adder #(4, 3, 0, 1, 5, 0, 1) op_766 (v628[3:0], v626[2:0], v766[4:0]); // 3.0
    wire [4:0] v767; shift_adder #(4, 2, 1, 1, 5, 2, 1) op_767 (v629[3:0], v413[1:0], v767[4:0]); // 3.0
    wire [4:0] v768; shift_adder #(5, 3, 1, 1, 5, 1, 0) op_768 (v630[4:0], v631[2:0], v768[4:0]); // 3.0
    wire [4:0] v769; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_769 (v632[2:0], v633[3:0], v769[4:0]); // 3.0
    wire [3:0] v770; shift_adder #(3, 3, 1, 1, 4, 0, 1) op_770 (v634[2:0], v623[2:0], v770[3:0]); // 3.0
    wire [2:0] v771; shift_adder #(2, 2, 1, 1, 3, 0, 1) op_771 (v636[1:0], v434[1:0], v771[2:0]); // 3.0
    wire [2:0] v772; shift_adder #(1, 3, 0, 1, 3, 0, 0) op_772 (v230[0:0], v637[2:0], v772[2:0]); // 3.0
    wire [2:0] v773; shift_adder #(1, 3, 0, 1, 3, 0, 1) op_773 (v233[0:0], v639[2:0], v773[2:0]); // 3.0
    wire [4:0] v774; shift_adder #(5, 2, 1, 0, 5, 1, 1) op_774 (v640[4:0], v441[1:0], v774[4:0]); // 3.0
    wire [4:0] v775; shift_adder #(4, 3, 0, 1, 5, 1, 1) op_775 (v641[3:0], v642[2:0], v775[4:0]); // 3.0
    wire [4:0] v776; shift_adder #(5, 3, 1, 1, 5, 2, 1) op_776 (v643[4:0], v447[2:0], v776[4:0]); // 3.0
    wire [3:0] v777; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_777 (v637[2:0], v645[2:0], v777[3:0]); // 3.0
    wire [4:0] v778; shift_adder #(3, 3, 1, 0, 5, -1, 0) op_778 (v647[2:0], v648[2:0], v778[4:0]); // 3.0
    wire [4:0] v779; shift_adder #(4, 3, 0, 1, 5, 0, 1) op_779 (v649[3:0], v647[2:0], v779[4:0]); // 3.0
    wire [4:0] v780; shift_adder #(4, 2, 1, 1, 5, 2, 1) op_780 (v650[3:0], v438[1:0], v780[4:0]); // 3.0
    wire [3:0] v781; shift_adder #(3, 3, 1, 1, 4, 0, 1) op_781 (v651[2:0], v642[2:0], v781[3:0]); // 3.0
    wire [4:0] v782; shift_adder #(5, 3, 1, 1, 5, 1, 0) op_782 (v653[4:0], v654[2:0], v782[4:0]); // 3.0
    wire [4:0] v783; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_783 (v655[2:0], v656[3:0], v783[4:0]); // 3.0
    wire [4:0] v784; shift_adder #(2, 5, 1, 1, 5, 0, 0) op_784 (v657[1:0], v658[4:0], v784[4:0]); // 3.0
    wire [2:0] v785; shift_adder #(1, 2, 0, 1, 3, 0, 0) op_785 (v212[0:0], v659[1:0], v785[2:0]); // 3.0
    wire [3:0] v786; shift_adder #(2, 4, 0, 1, 4, 0, 0) op_786 (v462[1:0], v660[3:0], v786[3:0]); // 3.0
    wire [4:0] v787; shift_adder #(4, 3, 1, 1, 5, -1, 1) op_787 (v662[3:0], v663[2:0], v787[4:0]); // 3.0
    wire [2:0] v788; shift_adder #(1, 2, 0, 1, 3, 0, 1) op_788 (v218[0:0], v659[1:0], v788[2:0]); // 3.0
    wire [4:0] v789; shift_adder #(5, 2, 1, 1, 5, 2, 1) op_789 (v664[4:0], v458[1:0], v789[4:0]); // 3.0
    wire [4:0] v790; shift_adder #(3, 3, 0, 0, 5, 1, 0) op_790 (v665[2:0], v469[2:0], v790[4:0]); // 3.0
    wire [3:0] v791; shift_adder #(3, 2, 1, 0, 4, 0, 1) op_791 (v667[2:0], v472[1:0], v791[3:0]); // 3.0
    wire [4:0] v792; shift_adder #(4, 2, 0, 0, 5, 1, 1) op_792 (v669[3:0], v461[1:0], v792[4:0]); // 3.0
    wire [5:0] v793; shift_adder #(5, 4, 1, 1, 6, 1, 1) op_793 (v670[4:0], v475[3:0], v793[5:0]); // 4.0
    wire [3:0] v794; shift_adder #(1, 3, 0, 1, 4, 0, 0) op_794 (v74[0:0], v671[2:0], v794[3:0]); // 4.0
    wire [6:0] v795; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_795 (v672[4:0], v673[4:0], v795[6:0]); // 4.0
    wire [6:0] v796; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_796 (v674[4:0], v675[4:0], v796[6:0]); // 4.0
    wire [3:0] v797; shift_adder #(1, 3, 0, 1, 4, 0, 0) op_797 (v131[0:0], v676[2:0], v797[3:0]); // 4.0
    wire [3:0] v798; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_798 (v677[2:0], v676[2:0], v798[3:0]); // 4.0
    wire [4:0] v799; shift_adder #(5, 3, 1, 1, 5, 0, 0) op_799 (v485[4:0], v678[2:0], v799[4:0]); // 4.0
    wire [4:0] v800; shift_adder #(5, 3, 1, 1, 5, 0, 1) op_800 (v679[4:0], v680[2:0], v800[4:0]); // 4.0
    wire [7:0] v801; shift_adder #(5, 4, 1, 0, 8, -3, 1) op_801 (v800[4:0], 4'b1001, v801[7:0]); // 4.0
    wire [6:0] v802; assign v802[6:0] = v801[6:0] & {7{~v801[7]}}; // 4.0
    wire [6:0] v803; shift_adder #(7, 4, 0, 0, 7, 0, 0) op_803 (v802[6:0], 4'b1000, v803[6:0]); // 4.0
    wire [2:0] v804; assign v804[2:0] = v803[6:4]; // 4.0
    wire [4:0] v805; shift_adder #(4, 3, 1, 1, 5, 1, 1) op_805 (v681[3:0], v491[2:0], v805[4:0]); // 4.0
    wire [3:0] v806; shift_adder #(1, 3, 0, 1, 4, 0, 0) op_806 (v80[0:0], v680[2:0], v806[3:0]); // 4.0
    wire [6:0] v807; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_807 (v684[4:0], v685[4:0], v807[6:0]); // 4.0
    wire [8:0] v808; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_808 (v807[6:0], 4'b1001, v808[8:0]); // 4.0
    wire [7:0] v809; assign v809[7:0] = v808[7:0] & {8{~v808[8]}}; // 4.0
    wire [7:0] v810; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_810 (v809[7:0], 4'b1000, v810[7:0]); // 4.0
    wire [3:0] v811; assign v811[3:0] = v810[7:4]; // 4.0
    wire [5:0] v812; shift_adder #(5, 3, 1, 1, 6, 1, 1) op_812 (v687[4:0], v491[2:0], v812[5:0]); // 4.0
    wire [3:0] v813; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_813 (v688[2:0], v671[2:0], v813[3:0]); // 4.0
    wire [4:0] v814; shift_adder #(5, 3, 1, 1, 5, 0, 0) op_814 (v503[4:0], v689[2:0], v814[4:0]); // 4.0
    wire [4:0] v815; shift_adder #(4, 4, 1, 1, 5, 0, 1) op_815 (v690[3:0], v506[3:0], v815[4:0]); // 4.0
    wire [8:0] v816; shift_adder #(5, 1, 1, 0, 9, -4, 0) op_816 (v815[4:0], 1'b1, v816[8:0]); // 4.0
    wire [6:0] v817; assign v817[6:0] = v816[6:0] & {7{~v816[8]}}; // 4.0
    wire [6:0] v818; shift_adder #(7, 5, 0, 0, 7, 0, 0) op_818 (v817[6:0], 5'b10000, v818[6:0]); // 4.0
    wire [1:0] v819; assign v819[1:0] = v818[6:5]; // 4.0
    wire [5:0] v820; shift_adder #(5, 3, 1, 1, 6, 1, 1) op_820 (v692[4:0], v510[2:0], v820[5:0]); // 4.0
    wire [4:0] v821; shift_adder #(4, 3, 1, 1, 5, 1, 1) op_821 (v693[3:0], v510[2:0], v821[4:0]); // 4.0
    wire [5:0] v822; shift_adder #(5, 4, 1, 0, 6, 1, 1) op_822 (v696[4:0], v515[3:0], v822[5:0]); // 4.0
    wire [6:0] v823; shift_adder #(6, 2, 1, 0, 7, -1, 0) op_823 (v822[5:0], 2'b11, v823[6:0]); // 4.0
    wire [4:0] v824; assign v824[4:0] = v823[4:0] & {5{~v823[6]}}; // 4.0
    wire [4:0] v825; shift_adder #(5, 3, 0, 0, 5, 0, 0) op_825 (v824[4:0], 3'b100, v825[4:0]); // 4.0
    wire [1:0] v826; assign v826[1:0] = v825[4:3]; // 4.0
    wire [5:0] v827; shift_adder #(5, 4, 1, 1, 6, 1, 0) op_827 (v697[4:0], v698[3:0], v827[5:0]); // 4.0
    wire [7:0] v828; shift_adder #(6, 4, 1, 0, 8, -2, 1) op_828 (v827[5:0], 4'b1001, v828[7:0]); // 4.0
    wire [6:0] v829; assign v829[6:0] = v828[6:0] & {7{~v828[7]}}; // 4.0
    wire [6:0] v830; shift_adder #(7, 4, 0, 0, 7, 0, 0) op_830 (v829[6:0], 4'b1000, v830[6:0]); // 4.0
    wire [2:0] v831; assign v831[2:0] = v830[6:4]; // 4.0
    wire [6:0] v832; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_832 (v699[4:0], v700[4:0], v832[6:0]); // 4.0
    wire [8:0] v833; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_833 (v832[6:0], 4'b1001, v833[8:0]); // 4.0
    wire [7:0] v834; assign v834[7:0] = v833[7:0] & {8{~v833[8]}}; // 4.0
    wire [7:0] v835; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_835 (v834[7:0], 4'b1000, v835[7:0]); // 4.0
    wire [3:0] v836; assign v836[3:0] = v835[7:4]; // 4.0
    wire [4:0] v837; shift_adder #(4, 4, 1, 1, 5, 0, 1) op_837 (v701[3:0], v524[3:0], v837[4:0]); // 4.0
    wire [5:0] v838; shift_adder #(5, 3, 1, 1, 6, 1, 1) op_838 (v703[4:0], v528[2:0], v838[5:0]); // 4.0
    wire [4:0] v839; shift_adder #(4, 4, 1, 1, 5, 0, 1) op_839 (v704[3:0], v530[3:0], v839[4:0]); // 4.0
    wire [6:0] v840; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_840 (v705[4:0], v706[4:0], v840[6:0]); // 4.0
    wire [8:0] v841; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_841 (v840[6:0], 4'b1001, v841[8:0]); // 4.0
    wire [7:0] v842; assign v842[7:0] = v841[7:0] & {8{~v841[8]}}; // 4.0
    wire [7:0] v843; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_843 (v842[7:0], 4'b1000, v843[7:0]); // 4.0
    wire [3:0] v844; assign v844[3:0] = v843[7:4]; // 4.0
    wire [3:0] v845; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_845 (v707[2:0], v708[2:0], v845[3:0]); // 4.0
    wire [4:0] v846; shift_adder #(5, 3, 1, 1, 5, 0, 0) op_846 (v537[4:0], v709[2:0], v846[4:0]); // 4.0
    wire [4:0] v847; shift_adder #(4, 3, 1, 1, 5, 1, 1) op_847 (v710[3:0], v528[2:0], v847[4:0]); // 4.0
    wire [4:0] v848; shift_adder #(4, 4, 1, 1, 5, 0, 1) op_848 (v712[3:0], v543[3:0], v848[4:0]); // 4.0
    wire [5:0] v849; shift_adder #(5, 4, 1, 1, 6, 1, 1) op_849 (v713[4:0], v545[3:0], v849[5:0]); // 4.0
    wire [5:0] v850; shift_adder #(5, 4, 1, 1, 6, 1, 1) op_850 (v714[4:0], v547[3:0], v850[5:0]); // 4.0
    wire [3:0] v851; shift_adder #(1, 3, 0, 1, 4, 0, 0) op_851 (v98[0:0], v708[2:0], v851[3:0]); // 4.0
    wire [3:0] v852; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_852 (v715[2:0], v716[2:0], v852[3:0]); // 4.0
    wire [4:0] v853; shift_adder #(5, 3, 1, 1, 5, 0, 0) op_853 (v550[4:0], v717[2:0], v853[4:0]); // 4.0
    wire [4:0] v854; shift_adder #(4, 4, 1, 1, 5, 0, 1) op_854 (v718[3:0], v554[3:0], v854[4:0]); // 4.0
    wire [4:0] v855; shift_adder #(4, 3, 1, 1, 5, 1, 1) op_855 (v719[3:0], v556[2:0], v855[4:0]); // 4.0
    wire [6:0] v856; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_856 (v721[4:0], v722[4:0], v856[6:0]); // 4.0
    wire [5:0] v857; shift_adder #(5, 4, 1, 1, 6, 1, 1) op_857 (v723[4:0], v562[3:0], v857[5:0]); // 4.0
    wire [3:0] v858; shift_adder #(1, 3, 0, 1, 4, 0, 0) op_858 (v89[0:0], v716[2:0], v858[3:0]); // 4.0
    wire [6:0] v859; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_859 (v724[4:0], v725[4:0], v859[6:0]); // 4.0
    wire [5:0] v860; shift_adder #(5, 3, 1, 1, 6, 1, 1) op_860 (v727[4:0], v556[2:0], v860[5:0]); // 4.0
    wire [6:0] v861; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_861 (v728[4:0], v729[4:0], v861[6:0]); // 4.0
    wire [8:0] v862; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_862 (v861[6:0], 4'b1001, v862[8:0]); // 4.0
    wire [7:0] v863; assign v863[7:0] = v862[7:0] & {8{~v862[8]}}; // 4.0
    wire [7:0] v864; shift_adder #(8, 3, 0, 0, 8, 0, 0) op_864 (v863[7:0], 3'b100, v864[7:0]); // 4.0
    wire [4:0] v865; assign v865[4:0] = v864[7:3]; // 4.0
    wire [5:0] v866; shift_adder #(3, 5, 1, 1, 6, -1, 0) op_866 (v730[2:0], v731[4:0], v866[5:0]); // 4.0
    wire [8:0] v867; shift_adder #(6, 2, 1, 0, 9, -3, 1) op_867 (v866[5:0], 2'b11, v867[8:0]); // 4.0
    wire [7:0] v868; assign v868[7:0] = v867[7:0] & {8{~v867[8]}}; // 4.0
    wire [7:0] v869; shift_adder #(8, 5, 0, 0, 8, 0, 0) op_869 (v868[7:0], 5'b10000, v869[7:0]); // 4.0
    wire [2:0] v870; assign v870[2:0] = v869[7:5]; // 4.0
    wire [3:0] v871; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_871 (v732[2:0], v733[2:0], v871[3:0]); // 4.0
    wire [4:0] v872; shift_adder #(5, 3, 1, 1, 5, 0, 0) op_872 (v575[4:0], v734[2:0], v872[4:0]); // 4.0
    wire [5:0] v873; shift_adder #(5, 4, 1, 1, 6, 1, 1) op_873 (v735[4:0], v578[3:0], v873[5:0]); // 4.0
    wire [3:0] v874; shift_adder #(1, 3, 0, 1, 4, 0, 0) op_874 (v140[0:0], v733[2:0], v874[3:0]); // 4.0
    wire [4:0] v875; shift_adder #(4, 3, 1, 1, 5, 1, 1) op_875 (v736[3:0], v580[2:0], v875[4:0]); // 4.0
    wire [5:0] v876; shift_adder #(5, 3, 1, 1, 6, 1, 1) op_876 (v739[4:0], v580[2:0], v876[5:0]); // 4.0
    wire [6:0] v877; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_877 (v740[4:0], v741[4:0], v877[6:0]); // 4.0
    wire [6:0] v878; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_878 (v742[4:0], v743[4:0], v878[6:0]); // 4.0
    wire [8:0] v879; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_879 (v878[6:0], 4'b1001, v879[8:0]); // 4.0
    wire [7:0] v880; assign v880[7:0] = v879[7:0] & {8{~v879[8]}}; // 4.0
    wire [7:0] v881; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_881 (v880[7:0], 4'b1000, v881[7:0]); // 4.0
    wire [3:0] v882; assign v882[3:0] = v881[7:4]; // 4.0
    wire [3:0] v883; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_883 (v744[2:0], v745[2:0], v883[3:0]); // 4.0
    wire [4:0] v884; shift_adder #(5, 3, 1, 1, 5, 0, 0) op_884 (v594[4:0], v746[2:0], v884[4:0]); // 4.0
    wire [5:0] v885; shift_adder #(5, 4, 1, 1, 6, 1, 1) op_885 (v747[4:0], v597[3:0], v885[5:0]); // 4.0
    wire [3:0] v886; shift_adder #(1, 3, 0, 1, 4, 0, 0) op_886 (v164[0:0], v745[2:0], v886[3:0]); // 4.0
    wire [6:0] v887; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_887 (v748[4:0], v749[4:0], v887[6:0]); // 4.0
    wire [4:0] v888; shift_adder #(4, 3, 1, 1, 5, 1, 1) op_888 (v750[3:0], v602[2:0], v888[4:0]); // 4.0
    wire [5:0] v889; shift_adder #(5, 3, 1, 1, 6, 1, 1) op_889 (v753[4:0], v602[2:0], v889[5:0]); // 4.0
    wire [6:0] v890; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_890 (v754[4:0], v755[4:0], v890[6:0]); // 4.0
    wire [8:0] v891; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_891 (v890[6:0], 4'b1001, v891[8:0]); // 4.0
    wire [7:0] v892; assign v892[7:0] = v891[7:0] & {8{~v891[8]}}; // 4.0
    wire [7:0] v893; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_893 (v892[7:0], 4'b1000, v893[7:0]); // 4.0
    wire [3:0] v894; assign v894[3:0] = v893[7:4]; // 4.0
    wire [4:0] v895; shift_adder #(4, 4, 1, 1, 5, 0, 1) op_895 (v756[3:0], v612[3:0], v895[4:0]); // 4.0
    wire [4:0] v896; shift_adder #(4, 4, 1, 1, 5, 0, 1) op_896 (v757[3:0], v614[3:0], v896[4:0]); // 4.0
    wire [3:0] v897; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_897 (v758[2:0], v759[2:0], v897[3:0]); // 4.0
    wire [4:0] v898; shift_adder #(5, 3, 1, 1, 5, 0, 0) op_898 (v617[4:0], v760[2:0], v898[4:0]); // 4.0
    wire [5:0] v899; shift_adder #(5, 4, 1, 1, 6, 1, 1) op_899 (v761[4:0], v620[3:0], v899[5:0]); // 4.0
    wire [3:0] v900; shift_adder #(1, 3, 0, 1, 4, 0, 0) op_900 (v182[0:0], v759[2:0], v900[3:0]); // 4.0
    wire [6:0] v901; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_901 (v762[4:0], v763[4:0], v901[6:0]); // 4.0
    wire [4:0] v902; shift_adder #(4, 3, 1, 1, 5, 1, 1) op_902 (v764[3:0], v625[2:0], v902[4:0]); // 4.0
    wire [5:0] v903; shift_adder #(5, 3, 1, 1, 6, 1, 1) op_903 (v767[4:0], v625[2:0], v903[5:0]); // 4.0
    wire [6:0] v904; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_904 (v768[4:0], v769[4:0], v904[6:0]); // 4.0
    wire [8:0] v905; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_905 (v904[6:0], 4'b1001, v905[8:0]); // 4.0
    wire [7:0] v906; assign v906[7:0] = v905[7:0] & {8{~v905[8]}}; // 4.0
    wire [7:0] v907; shift_adder #(8, 3, 0, 0, 8, 0, 0) op_907 (v906[7:0], 3'b100, v907[7:0]); // 4.0
    wire [4:0] v908; assign v908[4:0] = v907[7:3]; // 4.0
    wire [4:0] v909; shift_adder #(4, 4, 1, 1, 5, 0, 1) op_909 (v770[3:0], v635[3:0], v909[4:0]); // 4.0
    wire [3:0] v910; shift_adder #(3, 3, 1, 1, 4, 0, 0) op_910 (v771[2:0], v772[2:0], v910[3:0]); // 4.0
    wire [4:0] v911; shift_adder #(5, 3, 1, 1, 5, 0, 0) op_911 (v638[4:0], v773[2:0], v911[4:0]); // 4.0
    wire [6:0] v912; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_912 (v774[4:0], v775[4:0], v912[6:0]); // 4.0
    wire [3:0] v913; shift_adder #(1, 3, 0, 1, 4, 0, 0) op_913 (v200[0:0], v772[2:0], v913[3:0]); // 4.0
    wire [5:0] v914; shift_adder #(5, 4, 1, 1, 6, 1, 1) op_914 (v776[4:0], v644[3:0], v914[5:0]); // 4.0
    wire [4:0] v915; shift_adder #(4, 3, 1, 1, 5, 1, 1) op_915 (v777[3:0], v646[2:0], v915[4:0]); // 4.0
    wire [5:0] v916; shift_adder #(5, 3, 1, 1, 6, 1, 1) op_916 (v780[4:0], v646[2:0], v916[5:0]); // 4.0
    wire [4:0] v917; shift_adder #(4, 4, 1, 1, 5, 0, 1) op_917 (v781[3:0], v652[3:0], v917[4:0]); // 4.0
    wire [6:0] v918; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_918 (v782[4:0], v783[4:0], v918[6:0]); // 4.0
    wire [8:0] v919; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_919 (v918[6:0], 4'b1001, v919[8:0]); // 4.0
    wire [7:0] v920; assign v920[7:0] = v919[7:0] & {8{~v919[8]}}; // 4.0
    wire [7:0] v921; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_921 (v920[7:0], 4'b1000, v921[7:0]); // 4.0
    wire [3:0] v922; assign v922[3:0] = v921[7:4]; // 4.0
    wire [4:0] v923; shift_adder #(5, 3, 1, 1, 5, 0, 1) op_923 (v784[4:0], v785[2:0], v923[4:0]); // 4.0
    wire [6:0] v924; shift_adder #(5, 2, 1, 0, 7, -2, 0) op_924 (v923[4:0], 2'b11, v924[6:0]); // 4.0
    wire [5:0] v925; assign v925[5:0] = v924[5:0] & {6{~v924[6]}}; // 4.0
    wire [5:0] v926; shift_adder #(6, 2, 0, 0, 6, 0, 0) op_926 (v925[5:0], 2'b10, v926[5:0]); // 4.0
    wire [3:0] v927; assign v927[3:0] = v926[5:2]; // 4.0
    wire [4:0] v928; shift_adder #(4, 3, 1, 1, 5, 1, 1) op_928 (v786[3:0], v661[2:0], v928[4:0]); // 4.0
    wire [8:0] v929; shift_adder #(5, 2, 1, 0, 9, -4, 1) op_929 (v928[4:0], 2'b11, v929[8:0]); // 4.0
    wire [7:0] v930; assign v930[7:0] = v929[7:0] & {8{~v929[8]}}; // 4.0
    wire [7:0] v931; shift_adder #(8, 5, 0, 0, 8, 0, 0) op_931 (v930[7:0], 5'b10000, v931[7:0]); // 4.0
    wire [2:0] v932; assign v932[2:0] = v931[7:5]; // 4.0
    wire [4:0] v933; shift_adder #(5, 3, 1, 1, 5, 0, 1) op_933 (v787[4:0], v785[2:0], v933[4:0]); // 4.0
    wire [6:0] v934; shift_adder #(5, 3, 1, 0, 7, -2, 1) op_934 (v933[4:0], 3'b101, v934[6:0]); // 4.0
    wire [5:0] v935; assign v935[5:0] = v934[5:0] & {6{~v934[6]}}; // 4.0
    wire [5:0] v936; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_936 (v935[5:0], 3'b100, v936[5:0]); // 4.0
    wire [2:0] v937; assign v937[2:0] = v936[5:3]; // 4.0
    wire [2:0] v938; shift_adder #(1, 3, 0, 1, 3, -1, 1) op_938 (v212[0:0], v788[2:0], v938[2:0]); // 4.0
    wire [5:0] v939; shift_adder #(3, 5, 1, 1, 6, -2, 0) op_939 (v661[2:0], v789[4:0], v939[5:0]); // 4.0
    wire [4:0] v940; shift_adder #(4, 4, 1, 1, 5, 0, 0) op_940 (v666[3:0], v791[3:0], v940[4:0]); // 4.0
    wire [8:0] v941; shift_adder #(5, 1, 1, 0, 9, -4, 0) op_941 (v940[4:0], 1'b1, v941[8:0]); // 4.0
    wire [6:0] v942; assign v942[6:0] = v941[6:0] & {7{~v941[8]}}; // 4.0
    wire [6:0] v943; shift_adder #(7, 5, 0, 0, 7, 0, 0) op_943 (v942[6:0], 5'b10000, v943[6:0]); // 4.0
    wire [1:0] v944; assign v944[1:0] = v943[6:5]; // 4.0
    wire [5:0] v945; shift_adder #(3, 5, 0, 1, 6, -1, 0) op_945 (v668[2:0], v792[4:0], v945[5:0]); // 4.0
    wire [7:0] v946; shift_adder #(6, 4, 1, 0, 8, -2, 1) op_946 (v945[5:0], 4'b1001, v946[7:0]); // 4.0
    wire [6:0] v947; assign v947[6:0] = v946[6:0] & {7{~v946[7]}}; // 4.0
    wire [6:0] v948; shift_adder #(7, 4, 0, 0, 7, 0, 0) op_948 (v947[6:0], 4'b1000, v948[6:0]); // 4.0
    wire [2:0] v949; assign v949[2:0] = v948[6:4]; // 4.0
    wire [2:0] v950; shift_adder #(1, 4, 0, 1, 3, -1, 1) op_950 (v92[0:0], v794[3:0], v950[2:0]); // 5.0
    wire [2:0] v951; shift_adder #(1, 4, 0, 1, 3, -1, 1) op_951 (v128[0:0], v797[3:0], v951[2:0]); // 5.0
    wire [4:0] v952; shift_adder #(4, 5, 1, 1, 5, 0, 0) op_952 (v798[3:0], v799[4:0], v952[4:0]); // 5.0
    wire [6:0] v953; shift_adder #(5, 3, 1, 0, 7, -2, 1) op_953 (v952[4:0], 3'b101, v953[6:0]); // 5.0
    wire [5:0] v954; assign v954[5:0] = v953[5:0] & {6{~v953[6]}}; // 5.0
    wire [5:0] v955; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_955 (v954[5:0], 3'b100, v955[5:0]); // 5.0
    wire [2:0] v956; assign v956[2:0] = v955[5:3]; // 5.0
    wire [5:0] v957; shift_adder #(5, 5, 1, 1, 6, -1, 1) op_957 (v805[4:0], v682[4:0], v957[5:0]); // 5.0
    wire [6:0] v958; shift_adder #(6, 2, 1, 0, 7, -1, 0) op_958 (v957[5:0], 2'b11, v958[6:0]); // 5.0
    wire [5:0] v959; assign v959[5:0] = v958[5:0] & {6{~v958[6]}}; // 5.0
    wire [5:0] v960; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_960 (v959[5:0], 3'b100, v960[5:0]); // 5.0
    wire [2:0] v961; assign v961[2:0] = v960[5:3]; // 5.0
    wire [4:0] v962; shift_adder #(5, 4, 1, 1, 5, 0, 0) op_962 (v683[4:0], v806[3:0], v962[4:0]); // 5.0
    wire [6:0] v963; shift_adder #(5, 3, 1, 0, 7, -2, 1) op_963 (v962[4:0], 3'b101, v963[6:0]); // 5.0
    wire [5:0] v964; assign v964[5:0] = v963[5:0] & {6{~v963[6]}}; // 5.0
    wire [5:0] v965; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_965 (v964[5:0], 3'b100, v965[5:0]); // 5.0
    wire [2:0] v966; assign v966[2:0] = v965[5:3]; // 5.0
    wire [5:0] v967; shift_adder #(5, 6, 1, 1, 6, -1, 0) op_967 (v686[4:0], v812[5:0], v967[5:0]); // 5.0
    wire [8:0] v968; shift_adder #(6, 2, 1, 0, 9, -3, 1) op_968 (v967[5:0], 2'b11, v968[8:0]); // 5.0
    wire [7:0] v969; assign v969[7:0] = v968[7:0] & {8{~v968[8]}}; // 5.0
    wire [8:0] v970; shift_adder #(8, 5, 0, 0, 9, 0, 0) op_970 (v969[7:0], 5'b10000, v970[8:0]); // 5.0
    wire [3:0] v971; assign v971[3:0] = v970[8:5]; // 5.0
    wire [4:0] v972; shift_adder #(4, 5, 1, 1, 5, 0, 0) op_972 (v813[3:0], v814[4:0], v972[4:0]); // 5.0
    wire [6:0] v973; shift_adder #(5, 3, 1, 0, 7, -2, 1) op_973 (v972[4:0], 3'b101, v973[6:0]); // 5.0
    wire [5:0] v974; assign v974[5:0] = v973[5:0] & {6{~v973[6]}}; // 5.0
    wire [5:0] v975; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_975 (v974[5:0], 3'b100, v975[5:0]); // 5.0
    wire [2:0] v976; assign v976[2:0] = v975[5:3]; // 5.0
    wire [5:0] v977; shift_adder #(5, 6, 1, 1, 6, -1, 0) op_977 (v691[4:0], v820[5:0], v977[5:0]); // 5.0
    wire [8:0] v978; shift_adder #(6, 2, 1, 0, 9, -3, 1) op_978 (v977[5:0], 2'b11, v978[8:0]); // 5.0
    wire [7:0] v979; assign v979[7:0] = v978[7:0] & {8{~v978[8]}}; // 5.0
    wire [8:0] v980; shift_adder #(8, 5, 0, 0, 9, 0, 0) op_980 (v979[7:0], 5'b10000, v980[8:0]); // 5.0
    wire [3:0] v981; assign v981[3:0] = v980[8:5]; // 5.0
    wire [5:0] v982; shift_adder #(5, 5, 1, 1, 6, -1, 1) op_982 (v821[4:0], v694[4:0], v982[5:0]); // 5.0
    wire [6:0] v983; shift_adder #(6, 2, 1, 0, 7, -1, 0) op_983 (v982[5:0], 2'b11, v983[6:0]); // 5.0
    wire [5:0] v984; assign v984[5:0] = v983[5:0] & {6{~v983[6]}}; // 5.0
    wire [5:0] v985; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_985 (v984[5:0], 3'b100, v985[5:0]); // 5.0
    wire [2:0] v986; assign v986[2:0] = v985[5:3]; // 5.0
    wire [5:0] v987; shift_adder #(6, 4, 1, 1, 6, 1, 0) op_987 (v695[5:0], v806[3:0], v987[5:0]); // 5.0
    wire [5:0] v988; shift_adder #(6, 2, 1, 0, 6, 0, 1) op_988 (v987[5:0], 2'b10, v988[5:0]); // 5.0
    wire [4:0] v989; assign v989[4:0] = v988[4:0] & {5{~v988[5]}}; // 5.0
    wire [4:0] v990; shift_adder #(5, 2, 0, 0, 5, 0, 0) op_990 (v989[4:0], 2'b10, v990[4:0]); // 5.0
    wire [2:0] v991; assign v991[2:0] = v990[4:2]; // 5.0
    wire [3:0] v992; shift_adder #(2, 3, 0, 1, 4, 0, 0) op_992 (v826[1:0], v831[2:0], v992[3:0]); // 5.0
    wire [4:0] v993; shift_adder #(5, 3, 1, 1, 5, 1, 1) op_993 (v837[4:0], v689[2:0], v993[4:0]); // 5.0
    wire [8:0] v994; shift_adder #(5, 1, 1, 0, 9, -4, 0) op_994 (v993[4:0], 1'b1, v994[8:0]); // 5.0
    wire [7:0] v995; assign v995[7:0] = v994[7:0] & {8{~v994[8]}}; // 5.0
    wire [7:0] v996; shift_adder #(8, 5, 0, 0, 8, 0, 0) op_996 (v995[7:0], 5'b10000, v996[7:0]); // 5.0
    wire [2:0] v997; assign v997[2:0] = v996[7:5]; // 5.0
    wire [5:0] v998; shift_adder #(5, 6, 1, 1, 6, -1, 0) op_998 (v702[4:0], v838[5:0], v998[5:0]); // 5.0
    wire [8:0] v999; shift_adder #(6, 2, 1, 0, 9, -3, 1) op_999 (v998[5:0], 2'b11, v999[8:0]); // 5.0
    wire [7:0] v1000; assign v1000[7:0] = v999[7:0] & {8{~v999[8]}}; // 5.0
    wire [8:0] v1001; shift_adder #(8, 5, 0, 0, 9, 0, 0) op_1001 (v1000[7:0], 5'b10000, v1001[8:0]); // 5.0
    wire [3:0] v1002; assign v1002[3:0] = v1001[8:5]; // 5.0
    wire [4:0] v1003; shift_adder #(5, 3, 1, 1, 5, 1, 1) op_1003 (v839[4:0], v678[2:0], v1003[4:0]); // 5.0
    wire [8:0] v1004; shift_adder #(5, 1, 1, 0, 9, -4, 0) op_1004 (v1003[4:0], 1'b1, v1004[8:0]); // 5.0
    wire [7:0] v1005; assign v1005[7:0] = v1004[7:0] & {8{~v1004[8]}}; // 5.0
    wire [7:0] v1006; shift_adder #(8, 5, 0, 0, 8, 0, 0) op_1006 (v1005[7:0], 5'b10000, v1006[7:0]); // 5.0
    wire [2:0] v1007; assign v1007[2:0] = v1006[7:5]; // 5.0
    wire [4:0] v1008; shift_adder #(4, 5, 1, 1, 5, 0, 0) op_1008 (v845[3:0], v846[4:0], v1008[4:0]); // 5.0
    wire [6:0] v1009; shift_adder #(5, 3, 1, 0, 7, -2, 1) op_1009 (v1008[4:0], 3'b101, v1009[6:0]); // 5.0
    wire [5:0] v1010; assign v1010[5:0] = v1009[5:0] & {6{~v1009[6]}}; // 5.0
    wire [5:0] v1011; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_1011 (v1010[5:0], 3'b100, v1011[5:0]); // 5.0
    wire [2:0] v1012; assign v1012[2:0] = v1011[5:3]; // 5.0
    wire [5:0] v1013; shift_adder #(5, 5, 1, 1, 6, -1, 1) op_1013 (v847[4:0], v711[4:0], v1013[5:0]); // 5.0
    wire [6:0] v1014; shift_adder #(6, 2, 1, 0, 7, -1, 0) op_1014 (v1013[5:0], 2'b11, v1014[6:0]); // 5.0
    wire [5:0] v1015; assign v1015[5:0] = v1014[5:0] & {6{~v1014[6]}}; // 5.0
    wire [5:0] v1016; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_1016 (v1015[5:0], 3'b100, v1016[5:0]); // 5.0
    wire [2:0] v1017; assign v1017[2:0] = v1016[5:3]; // 5.0
    wire [4:0] v1018; shift_adder #(5, 3, 1, 1, 5, 1, 1) op_1018 (v848[4:0], v709[2:0], v1018[4:0]); // 5.0
    wire [8:0] v1019; shift_adder #(5, 1, 1, 0, 9, -4, 0) op_1019 (v1018[4:0], 1'b1, v1019[8:0]); // 5.0
    wire [7:0] v1020; assign v1020[7:0] = v1019[7:0] & {8{~v1019[8]}}; // 5.0
    wire [7:0] v1021; shift_adder #(8, 5, 0, 0, 8, 0, 0) op_1021 (v1020[7:0], 5'b10000, v1021[7:0]); // 5.0
    wire [2:0] v1022; assign v1022[2:0] = v1021[7:5]; // 5.0
    wire [2:0] v1023; shift_adder #(1, 4, 0, 1, 3, -1, 1) op_1023 (v83[0:0], v851[3:0], v1023[2:0]); // 5.0
    wire [4:0] v1024; shift_adder #(4, 5, 1, 1, 5, 0, 0) op_1024 (v852[3:0], v853[4:0], v1024[4:0]); // 5.0
    wire [6:0] v1025; shift_adder #(5, 3, 1, 0, 7, -2, 1) op_1025 (v1024[4:0], 3'b101, v1025[6:0]); // 5.0
    wire [5:0] v1026; assign v1026[5:0] = v1025[5:0] & {6{~v1025[6]}}; // 5.0
    wire [5:0] v1027; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_1027 (v1026[5:0], 3'b100, v1027[5:0]); // 5.0
    wire [2:0] v1028; assign v1028[2:0] = v1027[5:3]; // 5.0
    wire [4:0] v1029; shift_adder #(5, 3, 1, 1, 5, 1, 1) op_1029 (v854[4:0], v717[2:0], v1029[4:0]); // 5.0
    wire [8:0] v1030; shift_adder #(5, 1, 1, 0, 9, -4, 0) op_1030 (v1029[4:0], 1'b1, v1030[8:0]); // 5.0
    wire [7:0] v1031; assign v1031[7:0] = v1030[7:0] & {8{~v1030[8]}}; // 5.0
    wire [7:0] v1032; shift_adder #(8, 5, 0, 0, 8, 0, 0) op_1032 (v1031[7:0], 5'b10000, v1032[7:0]); // 5.0
    wire [2:0] v1033; assign v1033[2:0] = v1032[7:5]; // 5.0
    wire [5:0] v1034; shift_adder #(5, 5, 1, 1, 6, -1, 1) op_1034 (v855[4:0], v720[4:0], v1034[5:0]); // 5.0
    wire [6:0] v1035; shift_adder #(6, 2, 1, 0, 7, -1, 0) op_1035 (v1034[5:0], 2'b11, v1035[6:0]); // 5.0
    wire [5:0] v1036; assign v1036[5:0] = v1035[5:0] & {6{~v1035[6]}}; // 5.0
    wire [5:0] v1037; shift_adder #(6, 2, 0, 0, 6, 0, 0) op_1037 (v1036[5:0], 2'b10, v1037[5:0]); // 5.0
    wire [3:0] v1038; assign v1038[3:0] = v1037[5:2]; // 5.0
    wire [5:0] v1039; shift_adder #(4, 4, 1, 1, 6, -1, 1) op_1039 (v811[3:0], v836[3:0], v1039[5:0]); // 5.0
    wire [2:0] v1040; shift_adder #(1, 4, 0, 1, 3, -1, 1) op_1040 (v95[0:0], v858[3:0], v1040[2:0]); // 5.0
    wire [5:0] v1041; shift_adder #(5, 6, 1, 1, 6, -1, 0) op_1041 (v726[4:0], v860[5:0], v1041[5:0]); // 5.0
    wire [8:0] v1042; shift_adder #(6, 2, 1, 0, 9, -3, 1) op_1042 (v1041[5:0], 2'b11, v1042[8:0]); // 5.0
    wire [7:0] v1043; assign v1043[7:0] = v1042[7:0] & {8{~v1042[8]}}; // 5.0
    wire [8:0] v1044; shift_adder #(8, 5, 0, 0, 9, 0, 0) op_1044 (v1043[7:0], 5'b10000, v1044[8:0]); // 5.0
    wire [3:0] v1045; assign v1045[3:0] = v1044[8:5]; // 5.0
    wire [3:0] v1046; shift_adder #(3, 3, 0, 0, 4, -1, 0) op_1046 (v870[2:0], v804[2:0], v1046[3:0]); // 5.0
    wire [4:0] v1047; shift_adder #(3, 4, 1, 1, 5, -1, 1) op_1047 (v831[2:0], v811[3:0], v1047[4:0]); // 5.0
    wire [4:0] v1048; shift_adder #(2, 4, 0, 1, 5, 0, 0) op_1048 (v826[1:0], v811[3:0], v1048[4:0]); // 5.0
    wire [4:0] v1049; shift_adder #(4, 5, 1, 1, 5, 0, 0) op_1049 (v871[3:0], v872[4:0], v1049[4:0]); // 5.0
    wire [6:0] v1050; shift_adder #(5, 3, 1, 0, 7, -2, 1) op_1050 (v1049[4:0], 3'b101, v1050[6:0]); // 5.0
    wire [5:0] v1051; assign v1051[5:0] = v1050[5:0] & {6{~v1050[6]}}; // 5.0
    wire [5:0] v1052; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_1052 (v1051[5:0], 3'b100, v1052[5:0]); // 5.0
    wire [2:0] v1053; assign v1053[2:0] = v1052[5:3]; // 5.0
    wire [2:0] v1054; shift_adder #(1, 4, 0, 1, 3, -1, 1) op_1054 (v149[0:0], v874[3:0], v1054[2:0]); // 5.0
    wire [5:0] v1055; shift_adder #(5, 5, 1, 1, 6, -1, 1) op_1055 (v875[4:0], v737[4:0], v1055[5:0]); // 5.0
    wire [6:0] v1056; shift_adder #(6, 2, 1, 0, 7, -1, 0) op_1056 (v1055[5:0], 2'b11, v1056[6:0]); // 5.0
    wire [5:0] v1057; assign v1057[5:0] = v1056[5:0] & {6{~v1056[6]}}; // 5.0
    wire [5:0] v1058; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_1058 (v1057[5:0], 3'b100, v1058[5:0]); // 5.0
    wire [2:0] v1059; assign v1059[2:0] = v1058[5:3]; // 5.0
    wire [5:0] v1060; shift_adder #(5, 6, 1, 1, 6, -1, 0) op_1060 (v738[4:0], v876[5:0], v1060[5:0]); // 5.0
    wire [8:0] v1061; shift_adder #(6, 2, 1, 0, 9, -3, 1) op_1061 (v1060[5:0], 2'b11, v1061[8:0]); // 5.0
    wire [7:0] v1062; assign v1062[7:0] = v1061[7:0] & {8{~v1061[8]}}; // 5.0
    wire [8:0] v1063; shift_adder #(8, 5, 0, 0, 9, 0, 0) op_1063 (v1062[7:0], 5'b10000, v1063[8:0]); // 5.0
    wire [3:0] v1064; assign v1064[3:0] = v1063[8:5]; // 5.0
    wire [4:0] v1065; shift_adder #(4, 5, 1, 1, 5, 0, 0) op_1065 (v883[3:0], v884[4:0], v1065[4:0]); // 5.0
    wire [6:0] v1066; shift_adder #(5, 3, 1, 0, 7, -2, 1) op_1066 (v1065[4:0], 3'b101, v1066[6:0]); // 5.0
    wire [5:0] v1067; assign v1067[5:0] = v1066[5:0] & {6{~v1066[6]}}; // 5.0
    wire [5:0] v1068; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_1068 (v1067[5:0], 3'b100, v1068[5:0]); // 5.0
    wire [2:0] v1069; assign v1069[2:0] = v1068[5:3]; // 5.0
    wire [2:0] v1070; shift_adder #(1, 4, 0, 1, 3, -1, 1) op_1070 (v158[0:0], v886[3:0], v1070[2:0]); // 5.0
    wire [5:0] v1071; shift_adder #(5, 5, 1, 1, 6, -1, 1) op_1071 (v888[4:0], v751[4:0], v1071[5:0]); // 5.0
    wire [6:0] v1072; shift_adder #(6, 2, 1, 0, 7, -1, 0) op_1072 (v1071[5:0], 2'b11, v1072[6:0]); // 5.0
    wire [5:0] v1073; assign v1073[5:0] = v1072[5:0] & {6{~v1072[6]}}; // 5.0
    wire [5:0] v1074; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_1074 (v1073[5:0], 3'b100, v1074[5:0]); // 5.0
    wire [2:0] v1075; assign v1075[2:0] = v1074[5:3]; // 5.0
    wire [5:0] v1076; shift_adder #(5, 6, 1, 1, 6, -1, 0) op_1076 (v752[4:0], v889[5:0], v1076[5:0]); // 5.0
    wire [8:0] v1077; shift_adder #(6, 2, 1, 0, 9, -3, 1) op_1077 (v1076[5:0], 2'b11, v1077[8:0]); // 5.0
    wire [7:0] v1078; assign v1078[7:0] = v1077[7:0] & {8{~v1077[8]}}; // 5.0
    wire [8:0] v1079; shift_adder #(8, 5, 0, 0, 9, 0, 0) op_1079 (v1078[7:0], 5'b10000, v1079[8:0]); // 5.0
    wire [3:0] v1080; assign v1080[3:0] = v1079[8:5]; // 5.0
    wire [4:0] v1081; shift_adder #(5, 3, 1, 1, 5, 1, 1) op_1081 (v895[4:0], v746[2:0], v1081[4:0]); // 5.0
    wire [8:0] v1082; shift_adder #(5, 1, 1, 0, 9, -4, 0) op_1082 (v1081[4:0], 1'b1, v1082[8:0]); // 5.0
    wire [7:0] v1083; assign v1083[7:0] = v1082[7:0] & {8{~v1082[8]}}; // 5.0
    wire [7:0] v1084; shift_adder #(8, 5, 0, 0, 8, 0, 0) op_1084 (v1083[7:0], 5'b10000, v1084[7:0]); // 5.0
    wire [2:0] v1085; assign v1085[2:0] = v1084[7:5]; // 5.0
    wire [5:0] v1086; shift_adder #(4, 4, 1, 1, 6, -1, 1) op_1086 (v844[3:0], v882[3:0], v1086[5:0]); // 5.0
    wire [4:0] v1087; shift_adder #(5, 3, 1, 1, 5, 1, 1) op_1087 (v896[4:0], v734[2:0], v1087[4:0]); // 5.0
    wire [8:0] v1088; shift_adder #(5, 1, 1, 0, 9, -4, 0) op_1088 (v1087[4:0], 1'b1, v1088[8:0]); // 5.0
    wire [7:0] v1089; assign v1089[7:0] = v1088[7:0] & {8{~v1088[8]}}; // 5.0
    wire [7:0] v1090; shift_adder #(8, 5, 0, 0, 8, 0, 0) op_1090 (v1089[7:0], 5'b10000, v1090[7:0]); // 5.0
    wire [2:0] v1091; assign v1091[2:0] = v1090[7:5]; // 5.0
    wire [5:0] v1092; shift_adder #(4, 4, 1, 1, 6, -1, 1) op_1092 (v836[3:0], v844[3:0], v1092[5:0]); // 5.0
    wire [4:0] v1093; shift_adder #(4, 5, 1, 1, 5, 0, 0) op_1093 (v897[3:0], v898[4:0], v1093[4:0]); // 5.0
    wire [6:0] v1094; shift_adder #(5, 3, 1, 0, 7, -2, 1) op_1094 (v1093[4:0], 3'b101, v1094[6:0]); // 5.0
    wire [5:0] v1095; assign v1095[5:0] = v1094[5:0] & {6{~v1094[6]}}; // 5.0
    wire [5:0] v1096; shift_adder #(6, 2, 0, 0, 6, 0, 0) op_1096 (v1095[5:0], 2'b10, v1096[5:0]); // 5.0
    wire [3:0] v1097; assign v1097[3:0] = v1096[5:2]; // 5.0
    wire [2:0] v1098; shift_adder #(1, 4, 0, 1, 3, -1, 1) op_1098 (v176[0:0], v900[3:0], v1098[2:0]); // 5.0
    wire [5:0] v1099; shift_adder #(5, 5, 1, 1, 6, -1, 1) op_1099 (v902[4:0], v765[4:0], v1099[5:0]); // 5.0
    wire [6:0] v1100; shift_adder #(6, 2, 1, 0, 7, -1, 0) op_1100 (v1099[5:0], 2'b11, v1100[6:0]); // 5.0
    wire [5:0] v1101; assign v1101[5:0] = v1100[5:0] & {6{~v1100[6]}}; // 5.0
    wire [5:0] v1102; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_1102 (v1101[5:0], 3'b100, v1102[5:0]); // 5.0
    wire [2:0] v1103; assign v1103[2:0] = v1102[5:3]; // 5.0
    wire [5:0] v1104; shift_adder #(5, 6, 1, 1, 6, -1, 0) op_1104 (v766[4:0], v903[5:0], v1104[5:0]); // 5.0
    wire [8:0] v1105; shift_adder #(6, 2, 1, 0, 9, -3, 1) op_1105 (v1104[5:0], 2'b11, v1105[8:0]); // 5.0
    wire [7:0] v1106; assign v1106[7:0] = v1105[7:0] & {8{~v1105[8]}}; // 5.0
    wire [8:0] v1107; shift_adder #(8, 5, 0, 0, 9, 0, 0) op_1107 (v1106[7:0], 5'b10000, v1107[8:0]); // 5.0
    wire [3:0] v1108; assign v1108[3:0] = v1107[8:5]; // 5.0
    wire [4:0] v1109; shift_adder #(5, 3, 1, 1, 5, 1, 1) op_1109 (v909[4:0], v760[2:0], v1109[4:0]); // 5.0
    wire [8:0] v1110; shift_adder #(5, 1, 1, 0, 9, -4, 0) op_1110 (v1109[4:0], 1'b1, v1110[8:0]); // 5.0
    wire [7:0] v1111; assign v1111[7:0] = v1110[7:0] & {8{~v1110[8]}}; // 5.0
    wire [7:0] v1112; shift_adder #(8, 5, 0, 0, 8, 0, 0) op_1112 (v1111[7:0], 5'b10000, v1112[7:0]); // 5.0
    wire [2:0] v1113; assign v1113[2:0] = v1112[7:5]; // 5.0
    wire [5:0] v1114; shift_adder #(5, 4, 1, 1, 6, 0, 1) op_1114 (v865[4:0], v882[3:0], v1114[5:0]); // 5.0
    wire [4:0] v1115; shift_adder #(4, 5, 1, 1, 5, 0, 0) op_1115 (v910[3:0], v911[4:0], v1115[4:0]); // 5.0
    wire [6:0] v1116; shift_adder #(5, 3, 1, 0, 7, -2, 1) op_1116 (v1115[4:0], 3'b101, v1116[6:0]); // 5.0
    wire [5:0] v1117; assign v1117[5:0] = v1116[5:0] & {6{~v1116[6]}}; // 5.0
    wire [5:0] v1118; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_1118 (v1117[5:0], 3'b100, v1118[5:0]); // 5.0
    wire [2:0] v1119; assign v1119[2:0] = v1118[5:3]; // 5.0
    wire [2:0] v1120; shift_adder #(1, 4, 0, 1, 3, -1, 1) op_1120 (v194[0:0], v913[3:0], v1120[2:0]); // 5.0
    wire [5:0] v1121; shift_adder #(5, 5, 1, 1, 6, -1, 1) op_1121 (v915[4:0], v778[4:0], v1121[5:0]); // 5.0
    wire [6:0] v1122; shift_adder #(6, 2, 1, 0, 7, -1, 0) op_1122 (v1121[5:0], 2'b11, v1122[6:0]); // 5.0
    wire [5:0] v1123; assign v1123[5:0] = v1122[5:0] & {6{~v1122[6]}}; // 5.0
    wire [5:0] v1124; shift_adder #(6, 3, 0, 0, 6, 0, 0) op_1124 (v1123[5:0], 3'b100, v1124[5:0]); // 5.0
    wire [2:0] v1125; assign v1125[2:0] = v1124[5:3]; // 5.0
    wire [5:0] v1126; shift_adder #(5, 6, 1, 1, 6, -1, 0) op_1126 (v779[4:0], v916[5:0], v1126[5:0]); // 5.0
    wire [8:0] v1127; shift_adder #(6, 2, 1, 0, 9, -3, 1) op_1127 (v1126[5:0], 2'b11, v1127[8:0]); // 5.0
    wire [7:0] v1128; assign v1128[7:0] = v1127[7:0] & {8{~v1127[8]}}; // 5.0
    wire [8:0] v1129; shift_adder #(8, 5, 0, 0, 9, 0, 0) op_1129 (v1128[7:0], 5'b10000, v1129[8:0]); // 5.0
    wire [3:0] v1130; assign v1130[3:0] = v1129[8:5]; // 5.0
    wire [4:0] v1131; shift_adder #(5, 3, 1, 1, 5, 1, 1) op_1131 (v917[4:0], v773[2:0], v1131[4:0]); // 5.0
    wire [8:0] v1132; shift_adder #(5, 1, 1, 0, 9, -4, 0) op_1132 (v1131[4:0], 1'b1, v1132[8:0]); // 5.0
    wire [7:0] v1133; assign v1133[7:0] = v1132[7:0] & {8{~v1132[8]}}; // 5.0
    wire [7:0] v1134; shift_adder #(8, 5, 0, 0, 8, 0, 0) op_1134 (v1133[7:0], 5'b10000, v1134[7:0]); // 5.0
    wire [2:0] v1135; assign v1135[2:0] = v1134[7:5]; // 5.0
    wire [5:0] v1136; shift_adder #(4, 4, 1, 1, 6, -1, 1) op_1136 (v882[3:0], v894[3:0], v1136[5:0]); // 5.0
    wire [4:0] v1137; shift_adder #(4, 4, 1, 1, 5, 0, 0) op_1137 (v894[3:0], v922[3:0], v1137[4:0]); // 5.0
    wire [5:0] v1138; shift_adder #(3, 6, 1, 1, 6, -1, 0) op_1138 (v938[2:0], v939[5:0], v1138[5:0]); // 5.0
    wire [7:0] v1139; shift_adder #(6, 4, 1, 0, 8, -2, 1) op_1139 (v1138[5:0], 4'b1001, v1139[7:0]); // 5.0
    wire [6:0] v1140; assign v1140[6:0] = v1139[6:0] & {7{~v1139[7]}}; // 5.0
    wire [6:0] v1141; shift_adder #(7, 4, 0, 0, 7, 0, 0) op_1141 (v1140[6:0], 4'b1000, v1141[6:0]); // 5.0
    wire [2:0] v1142; assign v1142[2:0] = v1141[6:4]; // 5.0
    wire [5:0] v1143; shift_adder #(3, 5, 1, 0, 6, -1, 0) op_1143 (v938[2:0], v790[4:0], v1143[5:0]); // 5.0
    wire [5:0] v1144; shift_adder #(6, 2, 1, 0, 6, 0, 0) op_1144 (v1143[5:0], 2'b10, v1144[5:0]); // 5.0
    wire [5:0] v1144_neg; negative #(6, 6, 1) op_neg_1144 (v1144, v1144_neg);
    wire [2:0] v1145; assign v1145[2:0] = v1144_neg[2:0] & {3{~v1144_neg[5]}}; // 5.0
    wire [2:0] v1146; shift_adder #(3, 2, 0, 0, 3, 0, 0) op_1146 (v1145[2:0], 2'b10, v1146[2:0]); // 5.0
    wire [0:0] v1147; assign v1147[0:0] = v1146[2:2]; // 5.0
    wire [4:0] v1148; shift_adder #(4, 3, 1, 1, 5, 1, 1) op_1148 (v922[3:0], v932[2:0], v1148[4:0]); // 5.0
    wire [5:0] v1149; shift_adder #(4, 3, 0, 0, 6, 2, 1) op_1149 (v927[3:0], v949[2:0], v1149[5:0]); // 5.0
    wire [4:0] v1150; shift_adder #(3, 4, 0, 0, 5, 1, 0) op_1150 (v949[2:0], v927[3:0], v1150[4:0]); // 5.0
    wire [3:0] v1151; shift_adder #(2, 3, 0, 0, 4, -1, 0) op_1151 (v944[1:0], v949[2:0], v1151[3:0]); // 5.0
    wire [5:0] v1152; shift_adder #(5, 3, 1, 0, 6, 0, 1) op_1152 (v908[4:0], v949[2:0], v1152[5:0]); // 5.0
    wire [6:0] v1153; shift_adder #(5, 4, 1, 0, 7, -1, 1) op_1153 (v908[4:0], v927[3:0], v1153[6:0]); // 5.0
    wire [4:0] v1154; shift_adder #(3, 3, 1, 0, 5, 0, 0) op_1154 (v932[2:0], v949[2:0], v1154[4:0]); // 5.0
    wire [3:0] v1155; shift_adder #(2, 3, 0, 0, 4, 0, 1) op_1155 (v944[1:0], v937[2:0], v1155[3:0]); // 5.0
    wire [5:0] v1156; shift_adder #(4, 4, 1, 0, 6, 1, 1) op_1156 (v922[3:0], v927[3:0], v1156[5:0]); // 5.0
    wire [2:0] v1157; shift_adder #(2, 2, 0, 0, 3, 0, 0) op_1157 (v826[1:0], v819[1:0], v1157[2:0]); // 5.0
    wire [4:0] v1158; shift_adder #(3, 4, 0, 1, 5, 0, 1) op_1158 (v804[2:0], v811[3:0], v1158[4:0]); // 5.0
    wire [3:0] v1159; shift_adder #(3, 2, 1, 0, 4, 0, 1) op_1159 (v831[2:0], v826[1:0], v1159[3:0]); // 5.0
    wire [4:0] v1160; shift_adder #(3, 3, 0, 0, 5, 1, 1) op_1160 (v870[2:0], v804[2:0], v1160[4:0]); // 5.0
    wire [3:0] v1161; shift_adder #(2, 2, 0, 0, 4, -1, 0) op_1161 (v819[1:0], v826[1:0], v1161[3:0]); // 5.0
    wire [5:0] v1162; shift_adder #(4, 4, 1, 1, 6, -1, 1) op_1162 (v894[3:0], v922[3:0], v1162[5:0]); // 5.0
    wire [5:0] v1163; shift_adder #(6, 3, 1, 1, 6, 1, 1) op_1163 (v793[5:0], v950[2:0], v1163[5:0]); // 6.0
    wire [5:0] v1164; shift_adder #(6, 2, 1, 0, 6, 0, 1) op_1164 (v1163[5:0], 2'b10, v1164[5:0]); // 6.0
    wire [4:0] v1165; assign v1165[4:0] = v1164[4:0] & {5{~v1164[5]}}; // 6.0
    wire [4:0] v1166; shift_adder #(5, 1, 0, 0, 5, 0, 0) op_1166 (v1165[4:0], 1'b1, v1166[4:0]); // 6.0
    wire [3:0] v1167; assign v1167[3:0] = v1166[4:1]; // 6.0
    wire [6:0] v1168; shift_adder #(7, 3, 1, 1, 7, 1, 0) op_1168 (v795[6:0], v950[2:0], v1168[6:0]); // 6.0
    wire [8:0] v1169; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_1169 (v1168[6:0], 4'b1001, v1169[8:0]); // 6.0
    wire [7:0] v1170; assign v1170[7:0] = v1169[7:0] & {8{~v1169[8]}}; // 6.0
    wire [7:0] v1171; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_1171 (v1170[7:0], 4'b1000, v1171[7:0]); // 6.0
    wire [3:0] v1172; assign v1172[3:0] = v1171[7:4]; // 6.0
    wire [6:0] v1173; shift_adder #(7, 3, 1, 1, 7, 1, 0) op_1173 (v796[6:0], v951[2:0], v1173[6:0]); // 6.0
    wire [8:0] v1174; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_1174 (v1173[6:0], 4'b1001, v1174[8:0]); // 6.0
    wire [7:0] v1175; assign v1175[7:0] = v1174[7:0] & {8{~v1174[8]}}; // 6.0
    wire [7:0] v1176; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_1176 (v1175[7:0], 4'b1000, v1176[7:0]); // 6.0
    wire [3:0] v1177; assign v1177[3:0] = v1176[7:4]; // 6.0
    wire [3:0] v1178; shift_adder #(3, 3, 0, 0, 4, 0, 1) op_1178 (v804[2:0], v961[2:0], v1178[3:0]); // 6.0
    wire [4:0] v1179; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_1179 (v966[2:0], v811[3:0], v1179[4:0]); // 6.0
    wire [5:0] v1180; shift_adder #(4, 3, 1, 0, 6, 1, 0) op_1180 (v971[3:0], v976[2:0], v1180[5:0]); // 6.0
    wire [4:0] v1181; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1181 (v981[3:0], v986[2:0], v1181[4:0]); // 6.0
    wire [3:0] v1182; shift_adder #(3, 2, 0, 0, 4, 0, 1) op_1182 (v991[2:0], v819[1:0], v1182[3:0]); // 6.0
    wire [4:0] v1183; shift_adder #(4, 4, 1, 1, 5, 0, 0) op_1183 (v992[3:0], v981[3:0], v1183[4:0]); // 6.0
    wire [4:0] v1184; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1184 (v836[3:0], v976[2:0], v1184[4:0]); // 6.0
    wire [4:0] v1185; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1185 (v971[3:0], v986[2:0], v1185[4:0]); // 6.0
    wire [4:0] v1186; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1186 (v1002[3:0], v1007[2:0], v1186[4:0]); // 6.0
    wire [4:0] v1187; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1187 (v811[3:0], v961[2:0], v1187[4:0]); // 6.0
    wire [4:0] v1188; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1188 (v844[3:0], v1012[2:0], v1188[4:0]); // 6.0
    wire [4:0] v1189; shift_adder #(3, 3, 0, 0, 5, 1, 0) op_1189 (v1017[2:0], v1022[2:0], v1189[4:0]); // 6.0
    wire [5:0] v1190; shift_adder #(6, 3, 1, 1, 6, 1, 1) op_1190 (v849[5:0], v951[2:0], v1190[5:0]); // 6.0
    wire [5:0] v1191; shift_adder #(6, 2, 1, 0, 6, 0, 1) op_1191 (v1190[5:0], 2'b10, v1191[5:0]); // 6.0
    wire [4:0] v1192; assign v1192[4:0] = v1191[4:0] & {5{~v1191[5]}}; // 6.0
    wire [4:0] v1193; shift_adder #(5, 2, 0, 0, 5, 0, 0) op_1193 (v1192[4:0], 2'b10, v1193[4:0]); // 6.0
    wire [2:0] v1194; assign v1194[2:0] = v1193[4:2]; // 6.0
    wire [5:0] v1195; shift_adder #(6, 3, 1, 1, 6, 1, 1) op_1195 (v850[5:0], v1023[2:0], v1195[5:0]); // 6.0
    wire [5:0] v1196; shift_adder #(6, 2, 1, 0, 6, 0, 1) op_1196 (v1195[5:0], 2'b10, v1196[5:0]); // 6.0
    wire [4:0] v1197; assign v1197[4:0] = v1196[4:0] & {5{~v1196[5]}}; // 6.0
    wire [4:0] v1198; shift_adder #(5, 1, 0, 0, 5, 0, 0) op_1198 (v1197[4:0], 1'b1, v1198[4:0]); // 6.0
    wire [3:0] v1199; assign v1199[3:0] = v1198[4:1]; // 6.0
    wire [4:0] v1200; shift_adder #(3, 3, 0, 0, 5, -1, 0) op_1200 (v1017[2:0], v1028[2:0], v1200[4:0]); // 6.0
    wire [4:0] v1201; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1201 (v844[3:0], v986[2:0], v1201[4:0]); // 6.0
    wire [6:0] v1202; shift_adder #(7, 3, 1, 1, 7, 1, 0) op_1202 (v856[6:0], v1023[2:0], v1202[6:0]); // 6.0
    wire [8:0] v1203; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_1203 (v1202[6:0], 4'b1001, v1203[8:0]); // 6.0
    wire [7:0] v1204; assign v1204[7:0] = v1203[7:0] & {8{~v1203[8]}}; // 6.0
    wire [7:0] v1205; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_1205 (v1204[7:0], 4'b1000, v1205[7:0]); // 6.0
    wire [3:0] v1206; assign v1206[3:0] = v1205[7:4]; // 6.0
    wire [5:0] v1207; shift_adder #(4, 4, 1, 1, 6, 1, 1) op_1207 (v836[3:0], v1002[3:0], v1207[5:0]); // 6.0
    wire [5:0] v1208; shift_adder #(3, 4, 1, 1, 6, 1, 1) op_1208 (v831[2:0], v971[3:0], v1208[5:0]); // 6.0
    wire [4:0] v1209; shift_adder #(3, 3, 0, 0, 5, -1, 0) op_1209 (v986[2:0], v1012[2:0], v1209[4:0]); // 6.0
    wire [4:0] v1210; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1210 (v836[3:0], v961[2:0], v1210[4:0]); // 6.0
    wire [5:0] v1211; shift_adder #(4, 4, 1, 1, 6, 1, 1) op_1211 (v811[3:0], v981[3:0], v1211[5:0]); // 6.0
    wire [4:0] v1212; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_1212 (v956[2:0], v836[3:0], v1212[4:0]); // 6.0
    wire [5:0] v1213; shift_adder #(4, 3, 1, 0, 6, 1, 0) op_1213 (v981[3:0], v1012[2:0], v1213[5:0]); // 6.0
    wire [5:0] v1214; shift_adder #(3, 4, 0, 1, 6, -1, 0) op_1214 (v1007[2:0], v1002[3:0], v1214[5:0]); // 6.0
    wire [5:0] v1215; shift_adder #(3, 4, 0, 1, 6, 1, 1) op_1215 (v986[2:0], v844[3:0], v1215[5:0]); // 6.0
    wire [5:0] v1216; shift_adder #(4, 6, 1, 1, 6, 0, 0) op_1216 (v971[3:0], v1039[5:0], v1216[5:0]); // 6.0
    wire [4:0] v1217; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_1217 (v976[2:0], v844[3:0], v1217[4:0]); // 6.0
    wire [5:0] v1218; shift_adder #(4, 3, 1, 0, 6, 1, 0) op_1218 (v1002[3:0], v1028[2:0], v1218[5:0]); // 6.0
    wire [5:0] v1219; shift_adder #(6, 3, 1, 1, 6, 1, 1) op_1219 (v857[5:0], v1040[2:0], v1219[5:0]); // 6.0
    wire [5:0] v1220; shift_adder #(6, 2, 1, 0, 6, 0, 1) op_1220 (v1219[5:0], 2'b10, v1220[5:0]); // 6.0
    wire [4:0] v1221; assign v1221[4:0] = v1220[4:0] & {5{~v1220[5]}}; // 6.0
    wire [4:0] v1222; shift_adder #(5, 2, 0, 0, 5, 0, 0) op_1222 (v1221[4:0], 2'b10, v1222[4:0]); // 6.0
    wire [2:0] v1223; assign v1223[2:0] = v1222[4:2]; // 6.0
    wire [6:0] v1224; shift_adder #(7, 3, 1, 1, 7, 1, 0) op_1224 (v859[6:0], v1040[2:0], v1224[6:0]); // 6.0
    wire [8:0] v1225; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_1225 (v1224[6:0], 4'b1001, v1225[8:0]); // 6.0
    wire [7:0] v1226; assign v1226[7:0] = v1225[7:0] & {8{~v1225[8]}}; // 6.0
    wire [7:0] v1227; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_1227 (v1226[7:0], 4'b1000, v1227[7:0]); // 6.0
    wire [3:0] v1228; assign v1228[3:0] = v1227[7:4]; // 6.0
    wire [5:0] v1229; shift_adder #(3, 4, 0, 1, 6, -1, 0) op_1229 (v997[2:0], v1045[3:0], v1229[5:0]); // 6.0
    wire [4:0] v1230; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1230 (v1045[3:0], v997[2:0], v1230[4:0]); // 6.0
    wire [4:0] v1231; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1231 (v836[3:0], v986[2:0], v1231[4:0]); // 6.0
    wire [5:0] v1232; shift_adder #(5, 3, 1, 0, 6, 1, 0) op_1232 (v865[4:0], v1028[2:0], v1232[5:0]); // 6.0
    wire [5:0] v1233; shift_adder #(4, 3, 0, 0, 6, 2, 0) op_1233 (v1038[3:0], v1033[2:0], v1233[5:0]); // 6.0
    wire [5:0] v1234; shift_adder #(3, 4, 0, 1, 6, 1, 1) op_1234 (v961[2:0], v836[3:0], v1234[5:0]); // 6.0
    wire [6:0] v1235; shift_adder #(4, 5, 0, 1, 7, 1, 0) op_1235 (v1046[3:0], v1047[4:0], v1235[6:0]); // 6.0
    wire [3:0] v1236; shift_adder #(3, 3, 0, 0, 4, 0, 1) op_1236 (v976[2:0], v997[2:0], v1236[3:0]); // 6.0
    wire [6:0] v1237; shift_adder #(5, 3, 1, 0, 7, 2, 0) op_1237 (v1048[4:0], v961[2:0], v1237[6:0]); // 6.0
    wire [5:0] v1238; shift_adder #(6, 3, 1, 1, 6, 1, 1) op_1238 (v873[5:0], v1054[2:0], v1238[5:0]); // 6.0
    wire [5:0] v1239; shift_adder #(6, 2, 1, 0, 6, 0, 1) op_1239 (v1238[5:0], 2'b10, v1239[5:0]); // 6.0
    wire [4:0] v1240; assign v1240[4:0] = v1239[4:0] & {5{~v1239[5]}}; // 6.0
    wire [4:0] v1241; shift_adder #(5, 2, 0, 0, 5, 0, 0) op_1241 (v1240[4:0], 2'b10, v1241[4:0]); // 6.0
    wire [2:0] v1242; assign v1242[2:0] = v1241[4:2]; // 6.0
    wire [5:0] v1243; shift_adder #(3, 4, 0, 1, 6, -1, 0) op_1243 (v1022[2:0], v1064[3:0], v1243[5:0]); // 6.0
    wire [6:0] v1244; shift_adder #(7, 3, 1, 1, 7, 1, 0) op_1244 (v877[6:0], v1054[2:0], v1244[6:0]); // 6.0
    wire [8:0] v1245; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_1245 (v1244[6:0], 4'b1001, v1245[8:0]); // 6.0
    wire [7:0] v1246; assign v1246[7:0] = v1245[7:0] & {8{~v1245[8]}}; // 6.0
    wire [7:0] v1247; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_1247 (v1246[7:0], 4'b1000, v1247[7:0]); // 6.0
    wire [3:0] v1248; assign v1248[3:0] = v1247[7:4]; // 6.0
    wire [5:0] v1249; shift_adder #(4, 3, 1, 0, 6, 1, 0) op_1249 (v1045[3:0], v1012[2:0], v1249[5:0]); // 6.0
    wire [4:0] v1250; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_1250 (v1028[2:0], v882[3:0], v1250[4:0]); // 6.0
    wire [5:0] v1251; shift_adder #(4, 3, 1, 0, 6, 1, 0) op_1251 (v1064[3:0], v1069[2:0], v1251[5:0]); // 6.0
    wire [5:0] v1252; shift_adder #(6, 3, 1, 1, 6, 1, 1) op_1252 (v885[5:0], v1070[2:0], v1252[5:0]); // 6.0
    wire [5:0] v1253; shift_adder #(6, 2, 1, 0, 6, 0, 1) op_1253 (v1252[5:0], 2'b10, v1253[5:0]); // 6.0
    wire [4:0] v1254; assign v1254[4:0] = v1253[4:0] & {5{~v1253[5]}}; // 6.0
    wire [4:0] v1255; shift_adder #(5, 1, 0, 0, 5, 0, 0) op_1255 (v1254[4:0], 1'b1, v1255[4:0]); // 6.0
    wire [3:0] v1256; assign v1256[3:0] = v1255[4:1]; // 6.0
    wire [6:0] v1257; shift_adder #(7, 3, 1, 1, 7, 1, 0) op_1257 (v887[6:0], v1070[2:0], v1257[6:0]); // 6.0
    wire [8:0] v1258; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_1258 (v1257[6:0], 4'b1001, v1258[8:0]); // 6.0
    wire [7:0] v1259; assign v1259[7:0] = v1258[7:0] & {8{~v1258[8]}}; // 6.0
    wire [7:0] v1260; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_1260 (v1259[7:0], 4'b1000, v1260[7:0]); // 6.0
    wire [3:0] v1261; assign v1261[3:0] = v1260[7:4]; // 6.0
    wire [5:0] v1262; shift_adder #(3, 4, 0, 1, 6, -1, 0) op_1262 (v1033[2:0], v1080[3:0], v1262[5:0]); // 6.0
    wire [4:0] v1263; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1263 (v1080[3:0], v1033[2:0], v1263[4:0]); // 6.0
    wire [5:0] v1264; shift_adder #(5, 4, 1, 0, 6, 0, 0) op_1264 (v865[4:0], v1038[3:0], v1264[5:0]); // 6.0
    wire [4:0] v1265; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1265 (v894[3:0], v1069[2:0], v1265[4:0]); // 6.0
    wire [4:0] v1266; shift_adder #(3, 3, 0, 0, 5, 1, 0) op_1266 (v1075[2:0], v1085[2:0], v1266[4:0]); // 6.0
    wire [6:0] v1267; shift_adder #(4, 4, 0, 1, 7, 2, 0) op_1267 (v1038[3:0], v1002[3:0], v1267[6:0]); // 6.0
    wire [5:0] v1268; shift_adder #(4, 4, 1, 1, 6, 1, 1) op_1268 (v844[3:0], v1045[3:0], v1268[5:0]); // 6.0
    wire [4:0] v1269; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1269 (v1045[3:0], v1059[2:0], v1269[4:0]); // 6.0
    wire [4:0] v1270; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1270 (v1064[3:0], v1022[2:0], v1270[4:0]); // 6.0
    wire [4:0] v1271; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1271 (v844[3:0], v1017[2:0], v1271[4:0]); // 6.0
    wire [4:0] v1272; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1272 (v882[3:0], v1053[2:0], v1272[4:0]); // 6.0
    wire [5:0] v1273; shift_adder #(3, 5, 0, 1, 6, 0, 1) op_1273 (v1017[2:0], v865[4:0], v1273[5:0]); // 6.0
    wire [5:0] v1274; shift_adder #(4, 6, 1, 1, 6, 0, 0) op_1274 (v981[3:0], v1092[5:0], v1274[5:0]); // 6.0
    wire [4:0] v1275; shift_adder #(3, 3, 0, 0, 5, -1, 0) op_1275 (v1059[2:0], v1069[2:0], v1275[4:0]); // 6.0
    wire [5:0] v1276; shift_adder #(4, 4, 1, 0, 6, -1, 0) op_1276 (v882[3:0], v1038[3:0], v1276[5:0]); // 6.0
    wire [6:0] v1277; shift_adder #(5, 4, 1, 1, 7, 2, 1) op_1277 (v865[4:0], v1064[3:0], v1277[6:0]); // 6.0
    wire [3:0] v1278; shift_adder #(3, 3, 0, 0, 4, 0, 0) op_1278 (v1028[2:0], v1012[2:0], v1278[3:0]); // 6.0
    wire [4:0] v1279; shift_adder #(3, 4, 0, 0, 5, 1, 0) op_1279 (v1017[2:0], v1038[3:0], v1279[4:0]); // 6.0
    wire [3:0] v1280; shift_adder #(3, 3, 0, 0, 4, 0, 1) op_1280 (v1053[2:0], v1091[2:0], v1280[3:0]); // 6.0
    wire [4:0] v1281; shift_adder #(4, 4, 1, 1, 5, 0, 0) op_1281 (v1080[3:0], v1097[3:0], v1281[4:0]); // 6.0
    wire [4:0] v1282; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_1282 (v1053[2:0], v894[3:0], v1282[4:0]); // 6.0
    wire [5:0] v1283; shift_adder #(6, 3, 1, 1, 6, 1, 1) op_1283 (v899[5:0], v1098[2:0], v1283[5:0]); // 6.0
    wire [5:0] v1284; shift_adder #(6, 2, 1, 0, 6, 0, 1) op_1284 (v1283[5:0], 2'b10, v1284[5:0]); // 6.0
    wire [4:0] v1285; assign v1285[4:0] = v1284[4:0] & {5{~v1284[5]}}; // 6.0
    wire [4:0] v1286; shift_adder #(5, 2, 0, 0, 5, 0, 0) op_1286 (v1285[4:0], 2'b10, v1286[4:0]); // 6.0
    wire [2:0] v1287; assign v1287[2:0] = v1286[4:2]; // 6.0
    wire [6:0] v1288; shift_adder #(7, 3, 1, 1, 7, 1, 0) op_1288 (v901[6:0], v1098[2:0], v1288[6:0]); // 6.0
    wire [8:0] v1289; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_1289 (v1288[6:0], 4'b1001, v1289[8:0]); // 6.0
    wire [7:0] v1290; assign v1290[7:0] = v1289[7:0] & {8{~v1289[8]}}; // 6.0
    wire [7:0] v1291; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_1291 (v1290[7:0], 4'b1000, v1291[7:0]); // 6.0
    wire [3:0] v1292; assign v1292[3:0] = v1291[7:4]; // 6.0
    wire [5:0] v1293; shift_adder #(3, 4, 0, 1, 6, -1, 0) op_1293 (v1091[2:0], v1108[3:0], v1293[5:0]); // 6.0
    wire [5:0] v1294; shift_adder #(5, 4, 1, 1, 6, 0, 0) op_1294 (v908[4:0], v1097[3:0], v1294[5:0]); // 6.0
    wire [4:0] v1295; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1295 (v1108[3:0], v1091[2:0], v1295[4:0]); // 6.0
    wire [4:0] v1296; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1296 (v882[3:0], v1059[2:0], v1296[4:0]); // 6.0
    wire [4:0] v1297; shift_adder #(3, 3, 0, 0, 5, 1, 0) op_1297 (v1103[2:0], v1113[2:0], v1297[4:0]); // 6.0
    wire [5:0] v1298; shift_adder #(4, 4, 1, 1, 6, 1, 1) op_1298 (v882[3:0], v1080[3:0], v1298[5:0]); // 6.0
    wire [5:0] v1299; shift_adder #(4, 3, 1, 0, 6, 2, 0) op_1299 (v1097[3:0], v1075[2:0], v1299[5:0]); // 6.0
    wire [4:0] v1300; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1300 (v894[3:0], v1059[2:0], v1300[4:0]); // 6.0
    wire [5:0] v1301; shift_adder #(3, 4, 0, 1, 6, 1, 1) op_1301 (v1059[2:0], v894[3:0], v1301[5:0]); // 6.0
    wire [5:0] v1302; shift_adder #(4, 6, 1, 1, 6, 0, 0) op_1302 (v1045[3:0], v1114[5:0], v1302[5:0]); // 6.0
    wire [6:0] v1303; shift_adder #(7, 3, 1, 1, 7, 1, 0) op_1303 (v912[6:0], v1120[2:0], v1303[6:0]); // 6.0
    wire [8:0] v1304; shift_adder #(7, 4, 1, 0, 9, -2, 1) op_1304 (v1303[6:0], 4'b1001, v1304[8:0]); // 6.0
    wire [7:0] v1305; assign v1305[7:0] = v1304[7:0] & {8{~v1304[8]}}; // 6.0
    wire [7:0] v1306; shift_adder #(8, 4, 0, 0, 8, 0, 0) op_1306 (v1305[7:0], 4'b1000, v1306[7:0]); // 6.0
    wire [3:0] v1307; assign v1307[3:0] = v1306[7:4]; // 6.0
    wire [5:0] v1308; shift_adder #(6, 3, 1, 1, 6, 1, 1) op_1308 (v914[5:0], v1120[2:0], v1308[5:0]); // 6.0
    wire [5:0] v1309; shift_adder #(6, 2, 1, 0, 6, 0, 1) op_1309 (v1308[5:0], 2'b10, v1309[5:0]); // 6.0
    wire [4:0] v1310; assign v1310[4:0] = v1309[4:0] & {5{~v1309[5]}}; // 6.0
    wire [4:0] v1311; shift_adder #(5, 2, 0, 0, 5, 0, 0) op_1311 (v1310[4:0], 2'b10, v1311[4:0]); // 6.0
    wire [2:0] v1312; assign v1312[2:0] = v1311[4:2]; // 6.0
    wire [5:0] v1313; shift_adder #(3, 5, 0, 1, 6, -1, 0) op_1313 (v1069[2:0], v908[4:0], v1313[5:0]); // 6.0
    wire [5:0] v1314; shift_adder #(3, 4, 0, 1, 6, -1, 0) op_1314 (v1085[2:0], v1130[3:0], v1314[5:0]); // 6.0
    wire [5:0] v1315; shift_adder #(5, 3, 1, 0, 6, 1, 0) op_1315 (v908[4:0], v1075[2:0], v1315[5:0]); // 6.0
    wire [4:0] v1316; shift_adder #(3, 3, 0, 0, 5, -1, 0) op_1316 (v1103[2:0], v1119[2:0], v1316[4:0]); // 6.0
    wire [5:0] v1317; shift_adder #(4, 4, 1, 1, 6, 1, 1) op_1317 (v894[3:0], v1108[3:0], v1317[5:0]); // 6.0
    wire [5:0] v1318; shift_adder #(3, 4, 0, 1, 6, -2, 0) op_1318 (v1125[2:0], v1097[3:0], v1318[5:0]); // 6.0
    wire [5:0] v1319; shift_adder #(3, 5, 0, 1, 6, 0, 1) op_1319 (v1075[2:0], v908[4:0], v1319[5:0]); // 6.0
    wire [5:0] v1320; shift_adder #(4, 6, 1, 1, 6, 0, 0) op_1320 (v1064[3:0], v1136[5:0], v1320[5:0]); // 6.0
    wire [5:0] v1321; shift_adder #(5, 3, 1, 0, 6, 0, 1) op_1321 (v1137[4:0], v1085[2:0], v1321[5:0]); // 6.0
    wire [4:0] v1322; shift_adder #(3, 3, 0, 0, 5, 1, 0) op_1322 (v1125[2:0], v1135[2:0], v1322[4:0]); // 6.0
    wire [4:0] v1323; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_1323 (v1075[2:0], v1130[3:0], v1323[4:0]); // 6.0
    wire [4:0] v1324; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1324 (v922[3:0], v1119[2:0], v1324[4:0]); // 6.0
    wire [4:0] v1325; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1325 (v922[3:0], v1119[2:0], v1325[4:0]); // 6.0
    wire [4:0] v1326; shift_adder #(3, 3, 0, 1, 5, -1, 0) op_1326 (v1113[2:0], v932[2:0], v1326[4:0]); // 6.0
    wire [4:0] v1327; shift_adder #(1, 4, 0, 1, 5, 0, 0) op_1327 (v1147[0:0], v1130[3:0], v1327[4:0]); // 6.0
    wire [4:0] v1328; shift_adder #(2, 3, 0, 0, 5, 1, 0) op_1328 (v944[1:0], v1142[2:0], v1328[4:0]); // 6.0
    wire [3:0] v1329; shift_adder #(3, 3, 0, 0, 4, 0, 0) op_1329 (v1119[2:0], v949[2:0], v1329[3:0]); // 6.0
    wire [2:0] v1330; shift_adder #(1, 3, 0, 0, 3, -1, 0) op_1330 (v1147[0:0], v937[2:0], v1330[2:0]); // 6.0
    wire [4:0] v1331; shift_adder #(3, 3, 1, 0, 5, 1, 0) op_1331 (v932[2:0], v1135[2:0], v1331[4:0]); // 6.0
    wire [3:0] v1332; shift_adder #(3, 3, 0, 0, 4, 0, 0) op_1332 (v1142[2:0], v937[2:0], v1332[3:0]); // 6.0
    wire [4:0] v1333; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1333 (v922[3:0], v1135[2:0], v1333[4:0]); // 6.0
    wire [5:0] v1334; shift_adder #(3, 3, 0, 1, 6, -1, 1) op_1334 (v1125[2:0], v932[2:0], v1334[5:0]); // 6.0
    wire [5:0] v1335; shift_adder #(4, 5, 1, 1, 6, -1, 1) op_1335 (v1130[3:0], v1148[4:0], v1335[5:0]); // 6.0
    wire [5:0] v1336; shift_adder #(1, 6, 0, 1, 6, -2, 0) op_1336 (v1147[0:0], v1149[5:0], v1336[5:0]); // 6.0
    wire [3:0] v1337; shift_adder #(1, 3, 0, 0, 4, -1, 0) op_1337 (v1147[0:0], v1125[2:0], v1337[3:0]); // 6.0
    wire [4:0] v1338; shift_adder #(3, 4, 0, 0, 5, 0, 0) op_1338 (v1142[2:0], v1151[3:0], v1338[4:0]); // 6.0
    wire [6:0] v1339; shift_adder #(5, 4, 1, 1, 7, 2, 1) op_1339 (v908[4:0], v1130[3:0], v1339[6:0]); // 6.0
    wire [5:0] v1340; shift_adder #(4, 6, 1, 1, 6, 0, 0) op_1340 (v1108[3:0], v1152[5:0], v1340[5:0]); // 6.0
    wire [5:0] v1341; shift_adder #(3, 4, 0, 1, 6, 1, 1) op_1341 (v1125[2:0], v922[3:0], v1341[5:0]); // 6.0
    wire [2:0] v1342; shift_adder #(1, 3, 0, 0, 3, 0, 0) op_1342 (v1147[0:0], v1103[2:0], v1342[2:0]); // 6.0
    wire [7:0] v1343; shift_adder #(7, 5, 1, 1, 8, 2, 0) op_1343 (v1153[6:0], v1154[4:0], v1343[7:0]); // 6.0
    wire [4:0] v1344; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1344 (v1155[3:0], v1113[2:0], v1344[4:0]); // 6.0
    wire [4:0] v1345; shift_adder #(3, 3, 0, 0, 5, 2, 0) op_1345 (v1103[2:0], v1125[2:0], v1345[4:0]); // 6.0
    wire [6:0] v1346; shift_adder #(6, 4, 1, 1, 7, 1, 1) op_1346 (v1156[5:0], v1155[3:0], v1346[6:0]); // 6.0
    wire [5:0] v1347; shift_adder #(3, 5, 0, 1, 6, 1, 0) op_1347 (v1157[2:0], v1158[4:0], v1347[5:0]); // 6.0
    wire [3:0] v1348; shift_adder #(3, 3, 0, 0, 4, 0, 0) op_1348 (v870[2:0], v991[2:0], v1348[3:0]); // 6.0
    wire [4:0] v1349; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1349 (v971[3:0], v961[2:0], v1349[4:0]); // 6.0
    wire [4:0] v1350; shift_adder #(3, 4, 0, 1, 5, 1, 0) op_1350 (v870[2:0], v1159[3:0], v1350[4:0]); // 6.0
    wire [3:0] v1351; shift_adder #(3, 3, 0, 0, 4, 0, 0) op_1351 (v804[2:0], v966[2:0], v1351[3:0]); // 6.0
    wire [5:0] v1352; shift_adder #(4, 5, 1, 1, 6, -1, 1) op_1352 (v971[3:0], v1160[4:0], v1352[5:0]); // 6.0
    wire [4:0] v1353; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1353 (v811[3:0], v956[2:0], v1353[4:0]); // 6.0
    wire [3:0] v1354; shift_adder #(2, 3, 0, 0, 4, 0, 1) op_1354 (v826[1:0], v961[2:0], v1354[3:0]); // 6.0
    wire [5:0] v1355; shift_adder #(4, 3, 1, 0, 6, 1, 0) op_1355 (v1159[3:0], v956[2:0], v1355[5:0]); // 6.0
    wire [4:0] v1356; shift_adder #(3, 5, 0, 1, 5, 0, 0) op_1356 (v1007[2:0], v1160[4:0], v1356[4:0]); // 6.0
    wire [4:0] v1357; shift_adder #(3, 3, 0, 0, 5, 1, 0) op_1357 (v966[2:0], v991[2:0], v1357[4:0]); // 6.0
    wire [5:0] v1358; shift_adder #(3, 5, 0, 1, 6, 0, 1) op_1358 (v1103[2:0], v908[4:0], v1358[5:0]); // 6.0
    wire [5:0] v1359; shift_adder #(4, 6, 1, 1, 6, 0, 0) op_1359 (v1080[3:0], v1162[5:0], v1359[5:0]); // 6.0
    wire [5:0] v1360; shift_adder #(4, 4, 0, 1, 6, 1, 0) op_1360 (v1167[3:0], v1172[3:0], v1360[5:0]); // 7.0
    wire [4:0] v1361; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1361 (v1177[3:0], v956[2:0], v1361[4:0]); // 7.0
    wire [5:0] v1362; shift_adder #(4, 5, 1, 1, 6, 0, 0) op_1362 (v1178[3:0], v1179[4:0], v1362[5:0]); // 7.0
    wire [4:0] v1363; shift_adder #(2, 5, 0, 1, 5, -1, 0) op_1363 (v819[1:0], v1181[4:0], v1363[4:0]); // 7.0
    wire [4:0] v1364; shift_adder #(4, 4, 1, 1, 5, 0, 0) op_1364 (v1182[3:0], v1177[3:0], v1364[4:0]); // 7.0
    wire [6:0] v1365; shift_adder #(4, 5, 0, 1, 7, 1, 0) op_1365 (v1167[3:0], v1183[4:0], v1365[6:0]); // 7.0
    wire [6:0] v1366; shift_adder #(5, 5, 1, 1, 7, -1, 1) op_1366 (v1184[4:0], v1185[4:0], v1366[6:0]); // 7.0
    wire [4:0] v1367; shift_adder #(3, 4, 0, 1, 5, -1, 0) op_1367 (v997[2:0], v1178[3:0], v1367[4:0]); // 7.0
    wire [5:0] v1368; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_1368 (v1186[4:0], v1187[4:0], v1368[5:0]); // 7.0
    wire [5:0] v1369; shift_adder #(5, 5, 1, 0, 6, -1, 1) op_1369 (v1188[4:0], v1189[4:0], v1369[5:0]); // 7.0
    wire [5:0] v1370; shift_adder #(3, 4, 0, 1, 6, -1, 1) op_1370 (v1194[2:0], v981[3:0], v1370[5:0]); // 7.0
    wire [5:0] v1371; shift_adder #(4, 4, 1, 0, 6, -1, 0) op_1371 (v1172[3:0], v1199[3:0], v1371[5:0]); // 7.0
    wire [4:0] v1372; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1372 (v1177[3:0], v986[2:0], v1372[4:0]); // 7.0
    wire [4:0] v1373; shift_adder #(4, 3, 0, 0, 5, 1, 1) op_1373 (v1199[3:0], v1033[2:0], v1373[4:0]); // 7.0
    wire [5:0] v1374; shift_adder #(5, 4, 1, 0, 6, 1, 1) op_1374 (v1201[4:0], v1038[3:0], v1374[5:0]); // 7.0
    wire [4:0] v1375; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1375 (v1206[3:0], v1012[2:0], v1375[4:0]); // 7.0
    wire [4:0] v1376; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1376 (v1172[3:0], v1017[2:0], v1376[4:0]); // 7.0
    wire [4:0] v1377; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1377 (v1172[3:0], v956[2:0], v1377[4:0]); // 7.0
    wire [5:0] v1378; shift_adder #(5, 3, 1, 0, 6, 1, 1) op_1378 (v1184[4:0], v1194[2:0], v1378[5:0]); // 7.0
    wire [6:0] v1379; shift_adder #(6, 5, 1, 1, 7, 0, 0) op_1379 (v1208[5:0], v1179[4:0], v1379[6:0]); // 7.0
    wire [5:0] v1380; shift_adder #(3, 4, 0, 1, 6, 1, 0) op_1380 (v1007[2:0], v1177[3:0], v1380[5:0]); // 7.0
    wire [4:0] v1381; shift_adder #(4, 3, 0, 0, 5, 1, 1) op_1381 (v1167[3:0], v1022[2:0], v1381[4:0]); // 7.0
    wire [5:0] v1382; shift_adder #(5, 3, 1, 0, 6, 2, 1) op_1382 (v1210[4:0], v1017[2:0], v1382[5:0]); // 7.0
    wire [4:0] v1383; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1383 (v1172[3:0], v976[2:0], v1383[4:0]); // 7.0
    wire [6:0] v1384; shift_adder #(5, 6, 1, 1, 7, -1, 0) op_1384 (v1212[4:0], v1213[5:0], v1384[6:0]); // 7.0
    wire [5:0] v1385; shift_adder #(4, 4, 0, 1, 6, 1, 0) op_1385 (v1199[3:0], v1206[3:0], v1385[5:0]); // 7.0
    wire [5:0] v1386; shift_adder #(3, 6, 0, 1, 6, 0, 1) op_1386 (v1017[2:0], v1214[5:0], v1386[5:0]); // 7.0
    wire [5:0] v1387; shift_adder #(3, 4, 0, 1, 6, 1, 0) op_1387 (v997[2:0], v1172[3:0], v1387[5:0]); // 7.0
    wire [7:0] v1388; shift_adder #(6, 6, 1, 1, 8, 1, 0) op_1388 (v1215[5:0], v1216[5:0], v1388[7:0]); // 7.0
    wire [5:0] v1389; shift_adder #(4, 4, 0, 1, 6, 0, 0) op_1389 (v1167[3:0], v1177[3:0], v1389[5:0]); // 7.0
    wire [6:0] v1390; shift_adder #(5, 6, 1, 1, 7, -1, 0) op_1390 (v1217[4:0], v1218[5:0], v1390[6:0]); // 7.0
    wire [4:0] v1391; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_1391 (v1223[2:0], v1228[3:0], v1391[4:0]); // 7.0
    wire [6:0] v1392; shift_adder #(4, 6, 0, 1, 7, 1, 1) op_1392 (v1038[3:0], v1229[5:0], v1392[6:0]); // 7.0
    wire [5:0] v1393; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_1393 (v1230[4:0], v1231[4:0], v1393[5:0]); // 7.0
    wire [6:0] v1394; shift_adder #(6, 6, 1, 0, 7, -1, 1) op_1394 (v1232[5:0], v1233[5:0], v1394[6:0]); // 7.0
    wire [5:0] v1395; shift_adder #(4, 4, 0, 1, 6, 0, 1) op_1395 (v1167[3:0], v1002[3:0], v1395[5:0]); // 7.0
    wire [4:0] v1396; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1396 (v1206[3:0], v1223[2:0], v1396[4:0]); // 7.0
    wire [5:0] v1397; shift_adder #(5, 5, 1, 1, 6, 0, 1) op_1397 (v1188[4:0], v1212[4:0], v1397[5:0]); // 7.0
    wire [4:0] v1398; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1398 (v1206[3:0], v976[2:0], v1398[4:0]); // 7.0
    wire [5:0] v1399; shift_adder #(3, 6, 0, 1, 6, -1, 1) op_1399 (v1194[2:0], v1208[5:0], v1399[5:0]); // 7.0
    wire [7:0] v1400; shift_adder #(6, 7, 1, 1, 8, 0, 0) op_1400 (v1234[5:0], v1235[6:0], v1400[7:0]); // 7.0
    wire [5:0] v1401; shift_adder #(4, 3, 1, 0, 6, 2, 1) op_1401 (v1178[3:0], v986[2:0], v1401[5:0]); // 7.0
    wire [6:0] v1402; shift_adder #(4, 7, 1, 1, 7, -1, 0) op_1402 (v1236[3:0], v1237[6:0], v1402[6:0]); // 7.0
    wire [6:0] v1403; shift_adder #(6, 5, 1, 1, 7, 1, 1) op_1403 (v1232[5:0], v1217[4:0], v1403[6:0]); // 7.0
    wire [5:0] v1404; shift_adder #(3, 4, 0, 1, 6, 1, 0) op_1404 (v1022[2:0], v1206[3:0], v1404[5:0]); // 7.0
    wire [4:0] v1405; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1405 (v1228[3:0], v1012[2:0], v1405[4:0]); // 7.0
    wire [4:0] v1406; shift_adder #(3, 3, 0, 0, 5, -1, 0) op_1406 (v1053[2:0], v1242[2:0], v1406[4:0]); // 7.0
    wire [5:0] v1407; shift_adder #(3, 6, 0, 1, 6, 0, 1) op_1407 (v1059[2:0], v1243[5:0], v1407[5:0]); // 7.0
    wire [5:0] v1408; shift_adder #(4, 6, 1, 1, 6, 0, 0) op_1408 (v1248[3:0], v1249[5:0], v1408[5:0]); // 7.0
    wire [4:0] v1409; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1409 (v1228[3:0], v1028[2:0], v1409[4:0]); // 7.0
    wire [5:0] v1410; shift_adder #(4, 4, 1, 0, 6, -1, 1) op_1410 (v1206[3:0], v1038[3:0], v1410[5:0]); // 7.0
    wire [4:0] v1411; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1411 (v1248[3:0], v1053[2:0], v1411[4:0]); // 7.0
    wire [6:0] v1412; shift_adder #(5, 6, 1, 1, 7, -1, 0) op_1412 (v1250[4:0], v1251[5:0], v1412[6:0]); // 7.0
    wire [5:0] v1413; shift_adder #(4, 4, 0, 1, 6, 1, 0) op_1413 (v1256[3:0], v1261[3:0], v1413[5:0]); // 7.0
    wire [4:0] v1414; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1414 (v1228[3:0], v1059[2:0], v1414[4:0]); // 7.0
    wire [5:0] v1415; shift_adder #(3, 6, 0, 1, 6, 0, 1) op_1415 (v1075[2:0], v1262[5:0], v1415[5:0]); // 7.0
    wire [6:0] v1416; shift_adder #(5, 6, 1, 1, 7, -1, 0) op_1416 (v1263[4:0], v1264[5:0], v1416[6:0]); // 7.0
    wire [5:0] v1417; shift_adder #(5, 5, 1, 0, 6, -1, 1) op_1417 (v1265[4:0], v1266[4:0], v1417[5:0]); // 7.0
    wire [5:0] v1418; shift_adder #(3, 4, 0, 1, 6, -1, 1) op_1418 (v1223[2:0], v1064[3:0], v1418[5:0]); // 7.0
    wire [5:0] v1419; shift_adder #(4, 4, 1, 0, 6, -1, 0) op_1419 (v1248[3:0], v1256[3:0], v1419[5:0]); // 7.0
    wire [5:0] v1420; shift_adder #(3, 4, 0, 1, 6, 1, 0) op_1420 (v1033[2:0], v1228[3:0], v1420[5:0]); // 7.0
    wire [6:0] v1421; shift_adder #(3, 6, 0, 1, 7, -1, 1) op_1421 (v1223[2:0], v1268[5:0], v1421[6:0]); // 7.0
    wire [6:0] v1422; shift_adder #(6, 4, 1, 1, 7, -1, 0) op_1422 (v1086[5:0], v1206[3:0], v1422[6:0]); // 7.0
    wire [5:0] v1423; shift_adder #(4, 4, 0, 1, 6, 1, 0) op_1423 (v1199[3:0], v1228[3:0], v1423[5:0]); // 7.0
    wire [4:0] v1424; shift_adder #(3, 5, 0, 1, 5, 0, 0) op_1424 (v1242[2:0], v1270[4:0], v1424[4:0]); // 7.0
    wire [5:0] v1425; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_1425 (v1271[4:0], v1272[4:0], v1425[5:0]); // 7.0
    wire [7:0] v1426; shift_adder #(6, 6, 1, 1, 8, 1, 0) op_1426 (v1273[5:0], v1274[5:0], v1426[7:0]); // 7.0
    wire [5:0] v1427; shift_adder #(4, 4, 0, 1, 6, 0, 0) op_1427 (v1199[3:0], v1172[3:0], v1427[5:0]); // 7.0
    wire [3:0] v1428; shift_adder #(3, 3, 0, 0, 4, 0, 1) op_1428 (v1242[2:0], v1085[2:0], v1428[3:0]); // 7.0
    wire [6:0] v1429; shift_adder #(6, 3, 1, 0, 7, 3, 1) op_1429 (v1276[5:0], v1075[2:0], v1429[6:0]); // 7.0
    wire [5:0] v1430; shift_adder #(5, 5, 1, 1, 6, 0, 1) op_1430 (v1265[4:0], v1250[4:0], v1430[5:0]); // 7.0
    wire [5:0] v1431; shift_adder #(3, 4, 0, 1, 6, 1, 0) op_1431 (v1091[2:0], v1248[3:0], v1431[5:0]); // 7.0
    wire [4:0] v1432; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1432 (v1261[3:0], v1053[2:0], v1432[4:0]); // 7.0
    wire [5:0] v1433; shift_adder #(4, 5, 1, 1, 6, 0, 0) op_1433 (v1248[3:0], v1272[4:0], v1433[5:0]); // 7.0
    wire [4:0] v1434; shift_adder #(4, 3, 0, 0, 5, 1, 0) op_1434 (v1278[3:0], v1223[2:0], v1434[4:0]); // 7.0
    wire [5:0] v1435; shift_adder #(4, 3, 1, 0, 6, 1, 1) op_1435 (v1280[3:0], v1059[2:0], v1435[5:0]); // 7.0
    wire [4:0] v1436; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1436 (v1261[3:0], v1069[2:0], v1436[4:0]); // 7.0
    wire [6:0] v1437; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_1437 (v1281[4:0], v1282[4:0], v1437[6:0]); // 7.0
    wire [4:0] v1438; shift_adder #(3, 4, 0, 1, 5, 0, 0) op_1438 (v1287[2:0], v1292[3:0], v1438[4:0]); // 7.0
    wire [4:0] v1439; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1439 (v1248[3:0], v1075[2:0], v1439[4:0]); // 7.0
    wire [5:0] v1440; shift_adder #(3, 6, 0, 1, 6, 0, 1) op_1440 (v1103[2:0], v1293[5:0], v1440[5:0]); // 7.0
    wire [6:0] v1441; shift_adder #(6, 5, 1, 1, 7, 1, 0) op_1441 (v1294[5:0], v1295[4:0], v1441[6:0]); // 7.0
    wire [5:0] v1442; shift_adder #(5, 5, 1, 0, 6, -1, 1) op_1442 (v1296[4:0], v1297[4:0], v1442[5:0]); // 7.0
    wire [5:0] v1443; shift_adder #(3, 4, 0, 1, 6, -1, 1) op_1443 (v1242[2:0], v1080[3:0], v1443[5:0]); // 7.0
    wire [4:0] v1444; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1444 (v1261[3:0], v1287[2:0], v1444[4:0]); // 7.0
    wire [6:0] v1445; shift_adder #(6, 3, 1, 0, 7, 1, 1) op_1445 (v1294[5:0], v1069[2:0], v1445[6:0]); // 7.0
    wire [4:0] v1446; shift_adder #(4, 3, 0, 0, 5, 1, 1) op_1446 (v1256[3:0], v1113[2:0], v1446[4:0]); // 7.0
    wire [5:0] v1447; shift_adder #(3, 4, 0, 1, 6, 1, 0) op_1447 (v1085[2:0], v1261[3:0], v1447[5:0]); // 7.0
    wire [5:0] v1448; shift_adder #(4, 5, 1, 1, 6, 0, 1) op_1448 (v1292[3:0], v1282[4:0], v1448[5:0]); // 7.0
    wire [5:0] v1449; shift_adder #(5, 3, 1, 0, 6, 2, 1) op_1449 (v1300[4:0], v1103[2:0], v1449[5:0]); // 7.0
    wire [7:0] v1450; shift_adder #(6, 6, 1, 1, 8, 1, 0) op_1450 (v1301[5:0], v1302[5:0], v1450[7:0]); // 7.0
    wire [5:0] v1451; shift_adder #(3, 4, 0, 1, 6, -1, 0) op_1451 (v1242[2:0], v1228[3:0], v1451[5:0]); // 7.0
    wire [4:0] v1452; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1452 (v1261[3:0], v1103[2:0], v1452[4:0]); // 7.0
    wire [4:0] v1453; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1453 (v1292[3:0], v1119[2:0], v1453[4:0]); // 7.0
    wire [4:0] v1454; shift_adder #(4, 3, 1, 0, 5, 0, 0) op_1454 (v1108[3:0], v1312[2:0], v1454[4:0]); // 7.0
    wire [6:0] v1455; shift_adder #(4, 6, 1, 1, 7, 0, 0) op_1455 (v1097[3:0], v1313[5:0], v1455[6:0]); // 7.0
    wire [5:0] v1456; shift_adder #(3, 6, 0, 1, 6, 0, 1) op_1456 (v1125[2:0], v1314[5:0], v1456[5:0]); // 7.0
    wire [3:0] v1457; shift_adder #(3, 3, 0, 0, 4, 0, 1) op_1457 (v1287[2:0], v1135[2:0], v1457[3:0]); // 7.0
    wire [7:0] v1458; shift_adder #(6, 5, 1, 0, 8, 2, 0) op_1458 (v1315[5:0], v1316[4:0], v1458[7:0]); // 7.0
    wire [6:0] v1459; shift_adder #(6, 4, 1, 1, 7, 1, 0) op_1459 (v1318[5:0], v1292[3:0], v1459[6:0]); // 7.0
    wire [7:0] v1460; shift_adder #(6, 6, 1, 1, 8, 1, 0) op_1460 (v1319[5:0], v1320[5:0], v1460[7:0]); // 7.0
    wire [5:0] v1461; shift_adder #(4, 4, 0, 1, 6, 0, 0) op_1461 (v1256[3:0], v1248[3:0], v1461[5:0]); // 7.0
    wire [6:0] v1462; shift_adder #(6, 5, 1, 0, 7, -1, 1) op_1462 (v1321[5:0], v1322[4:0], v1462[6:0]); // 7.0
    wire [5:0] v1463; shift_adder #(3, 5, 0, 1, 6, 0, 0) op_1463 (v1312[2:0], v1323[4:0], v1463[5:0]); // 7.0
    wire [5:0] v1464; shift_adder #(4, 4, 0, 1, 6, 0, 1) op_1464 (v1256[3:0], v1108[3:0], v1464[5:0]); // 7.0
    wire [5:0] v1465; shift_adder #(3, 4, 0, 1, 6, 1, 0) op_1465 (v1113[2:0], v1292[3:0], v1465[5:0]); // 7.0
    wire [5:0] v1466; shift_adder #(5, 4, 1, 0, 6, 0, 0) op_1466 (v1324[4:0], v1307[3:0], v1466[5:0]); // 7.0
    wire [6:0] v1467; shift_adder #(4, 5, 1, 1, 7, 1, 0) op_1467 (v1097[3:0], v1325[4:0], v1467[6:0]); // 7.0
    wire [5:0] v1468; shift_adder #(4, 5, 0, 1, 6, 1, 1) op_1468 (v927[3:0], v1326[4:0], v1468[5:0]); // 7.0
    wire [4:0] v1469; shift_adder #(4, 3, 1, 0, 5, 0, 1) op_1469 (v1292[3:0], v1125[2:0], v1469[4:0]); // 7.0
    wire [4:0] v1470; shift_adder #(3, 5, 0, 1, 5, 0, 0) op_1470 (v1142[2:0], v1327[4:0], v1470[4:0]); // 7.0
    wire [5:0] v1471; shift_adder #(4, 4, 0, 0, 6, -1, 1) op_1471 (v1307[3:0], v927[3:0], v1471[5:0]); // 7.0
    wire [5:0] v1472; shift_adder #(5, 4, 0, 0, 6, -1, 0) op_1472 (v1328[4:0], v1329[3:0], v1472[5:0]); // 7.0
    wire [4:0] v1473; shift_adder #(3, 3, 0, 0, 5, 1, 0) op_1473 (v1330[2:0], v1135[2:0], v1473[4:0]); // 7.0
    wire [6:0] v1474; shift_adder #(5, 4, 1, 0, 7, 1, 0) op_1474 (v1331[4:0], v1329[3:0], v1474[6:0]); // 7.0
    wire [3:0] v1475; shift_adder #(3, 3, 0, 0, 4, 0, 0) op_1475 (v1142[2:0], v1312[2:0], v1475[3:0]); // 7.0
    wire [5:0] v1476; shift_adder #(5, 6, 1, 1, 6, -1, 0) op_1476 (v1333[4:0], v1334[5:0], v1476[5:0]); // 7.0
    wire [6:0] v1477; shift_adder #(5, 6, 0, 1, 7, 0, 0) op_1477 (v1328[4:0], v1335[5:0], v1477[6:0]); // 7.0
    wire [6:0] v1478; shift_adder #(6, 4, 1, 0, 7, 1, 0) op_1478 (v1336[5:0], v1307[3:0], v1478[6:0]); // 7.0
    wire [5:0] v1479; shift_adder #(5, 4, 0, 0, 6, 0, 0) op_1479 (v1150[4:0], v1337[3:0], v1479[5:0]); // 7.0
    wire [5:0] v1480; shift_adder #(5, 3, 0, 0, 6, 1, 1) op_1480 (v1338[4:0], v1312[2:0], v1480[5:0]); // 7.0
    wire [4:0] v1481; shift_adder #(3, 4, 0, 0, 5, 1, 0) op_1481 (v1135[2:0], v1307[3:0], v1481[4:0]); // 7.0
    wire [7:0] v1482; shift_adder #(3, 7, 0, 1, 8, -2, 1) op_1482 (v1312[2:0], v1339[6:0], v1482[7:0]); // 7.0
    wire [5:0] v1483; shift_adder #(4, 6, 1, 1, 6, 0, 0) op_1483 (v1292[3:0], v1341[5:0], v1483[5:0]); // 7.0
    wire [7:0] v1484; shift_adder #(3, 8, 0, 1, 8, -2, 0) op_1484 (v1342[2:0], v1343[7:0], v1484[7:0]); // 7.0
    wire [5:0] v1485; shift_adder #(3, 4, 0, 1, 6, -1, 1) op_1485 (v1287[2:0], v1130[3:0], v1485[5:0]); // 7.0
    wire [5:0] v1486; shift_adder #(5, 3, 0, 0, 6, 1, 1) op_1486 (v1345[4:0], v1119[2:0], v1486[5:0]); // 7.0
    wire [6:0] v1487; shift_adder #(6, 4, 1, 0, 7, 1, 0) op_1487 (v1347[5:0], v1348[3:0], v1487[6:0]); // 7.0
    wire [5:0] v1488; shift_adder #(3, 5, 1, 1, 6, 0, 0) op_1488 (v831[2:0], v1349[4:0], v1488[5:0]); // 7.0
    wire [4:0] v1489; shift_adder #(3, 3, 0, 0, 5, -1, 0) op_1489 (v956[2:0], v1194[2:0], v1489[4:0]); // 7.0
    wire [5:0] v1490; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_1490 (v1349[4:0], v1350[4:0], v1490[5:0]); // 7.0
    wire [5:0] v1491; shift_adder #(4, 4, 1, 0, 6, 1, 0) op_1491 (v1177[3:0], v1351[3:0], v1491[5:0]); // 7.0
    wire [6:0] v1492; shift_adder #(3, 6, 0, 1, 7, -1, 0) op_1492 (v1194[2:0], v1352[5:0], v1492[6:0]); // 7.0
    wire [4:0] v1493; shift_adder #(4, 3, 1, 0, 5, 1, 1) op_1493 (v1354[3:0], v1007[2:0], v1493[4:0]); // 7.0
    wire [6:0] v1494; shift_adder #(6, 4, 1, 0, 7, 1, 0) op_1494 (v1355[5:0], v1348[3:0], v1494[6:0]); // 7.0
    wire [5:0] v1495; shift_adder #(4, 3, 1, 0, 6, -1, 1) op_1495 (v1354[3:0], v1007[2:0], v1495[5:0]); // 7.0
    wire [4:0] v1496; shift_adder #(4, 4, 1, 0, 5, 0, 1) op_1496 (v1177[3:0], v1161[3:0], v1496[4:0]); // 7.0
    wire [6:0] v1497; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_1497 (v1353[4:0], v1356[4:0], v1497[6:0]); // 7.0
    wire [7:0] v1498; shift_adder #(6, 6, 1, 1, 8, 1, 0) op_1498 (v1358[5:0], v1359[5:0], v1498[7:0]); // 7.0
    wire [5:0] v1499; shift_adder #(3, 4, 0, 1, 6, -1, 0) op_1499 (v1287[2:0], v1261[3:0], v1499[5:0]); // 7.0
    wire [7:0] v1500; shift_adder #(6, 5, 1, 1, 8, 2, 0) op_1500 (v1360[5:0], v1361[4:0], v1500[7:0]); // 8.0
    wire [6:0] v1501; shift_adder #(6, 5, 1, 1, 7, 0, 0) op_1501 (v1180[5:0], v1363[4:0], v1501[6:0]); // 8.0
    wire [6:0] v1502; shift_adder #(5, 7, 1, 1, 7, -1, 0) op_1502 (v1364[4:0], v1365[6:0], v1502[6:0]); // 8.0
    wire [6:0] v1503; shift_adder #(7, 5, 1, 1, 7, 0, 1) op_1503 (v1366[6:0], v1367[4:0], v1503[6:0]); // 8.0
    wire [7:0] v1504; shift_adder #(6, 6, 1, 1, 8, -1, 0) op_1504 (v1368[5:0], v1369[5:0], v1504[7:0]); // 8.0
    wire [6:0] v1505; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_1505 (v1370[5:0], v1371[5:0], v1505[6:0]); // 8.0
    wire [6:0] v1506; shift_adder #(5, 5, 0, 1, 7, -1, 0) op_1506 (v1200[4:0], v1373[4:0], v1506[6:0]); // 8.0
    wire [6:0] v1507; shift_adder #(6, 5, 1, 1, 7, 1, 1) op_1507 (v1374[5:0], v1375[4:0], v1507[6:0]); // 8.0
    wire [6:0] v1508; shift_adder #(5, 6, 1, 1, 7, 0, 1) op_1508 (v1376[4:0], v1207[5:0], v1508[6:0]); // 8.0
    wire [6:0] v1509; shift_adder #(5, 6, 1, 1, 7, 0, 0) op_1509 (v1377[4:0], v1378[5:0], v1509[6:0]); // 8.0
    wire [5:0] v1510; shift_adder #(5, 5, 1, 1, 6, 0, 1) op_1510 (v1367[4:0], v1363[4:0], v1510[5:0]); // 8.0
    wire [7:0] v1511; shift_adder #(7, 6, 1, 1, 8, 1, 0) op_1511 (v1379[6:0], v1380[5:0], v1511[7:0]); // 8.0
    wire [6:0] v1512; shift_adder #(5, 5, 0, 1, 7, -1, 0) op_1512 (v1209[4:0], v1381[4:0], v1512[6:0]); // 8.0
    wire [6:0] v1513; shift_adder #(6, 5, 1, 1, 7, 1, 1) op_1513 (v1382[5:0], v1383[4:0], v1513[6:0]); // 8.0
    wire [6:0] v1514; shift_adder #(5, 6, 1, 1, 7, 0, 1) op_1514 (v1372[4:0], v1211[5:0], v1514[6:0]); // 8.0
    wire [7:0] v1515; shift_adder #(5, 7, 1, 1, 8, -1, 0) op_1515 (v1383[4:0], v1384[6:0], v1515[7:0]); // 8.0
    wire [7:0] v1516; shift_adder #(6, 5, 1, 1, 8, 2, 0) op_1516 (v1385[5:0], v1372[4:0], v1516[7:0]); // 8.0
    wire [6:0] v1517; shift_adder #(6, 6, 1, 1, 7, 0, 1) op_1517 (v1387[5:0], v1211[5:0], v1517[6:0]); // 8.0
    wire [6:0] v1518; shift_adder #(6, 6, 1, 1, 7, 1, 0) op_1518 (v1389[5:0], v1386[5:0], v1518[6:0]); // 8.0
    wire [7:0] v1519; shift_adder #(5, 7, 1, 1, 8, -1, 0) op_1519 (v1375[4:0], v1390[6:0], v1519[7:0]); // 8.0
    wire [6:0] v1520; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_1520 (v1391[4:0], v1376[4:0], v1520[6:0]); // 8.0
    wire [8:0] v1521; shift_adder #(6, 7, 1, 1, 9, -2, 0) op_1521 (v1393[5:0], v1394[6:0], v1521[8:0]); // 8.0
    wire [6:0] v1522; shift_adder #(6, 5, 1, 1, 7, 1, 0) op_1522 (v1395[5:0], v1396[4:0], v1522[6:0]); // 8.0
    wire [6:0] v1523; shift_adder #(6, 5, 1, 1, 7, 0, 1) op_1523 (v1397[5:0], v1381[4:0], v1523[6:0]); // 8.0
    wire [5:0] v1524; shift_adder #(5, 6, 1, 1, 6, 0, 0) op_1524 (v1398[4:0], v1386[5:0], v1524[5:0]); // 8.0
    wire [6:0] v1525; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_1525 (v1380[5:0], v1399[5:0], v1525[6:0]); // 8.0
    wire [7:0] v1526; shift_adder #(8, 5, 1, 1, 8, 1, 1) op_1526 (v1400[7:0], v1363[4:0], v1526[7:0]); // 8.0
    wire [6:0] v1527; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_1527 (v1401[5:0], v1399[5:0], v1527[6:0]); // 8.0
    wire [6:0] v1528; shift_adder #(7, 5, 1, 1, 7, 1, 1) op_1528 (v1402[6:0], v1361[4:0], v1528[6:0]); // 8.0
    wire [7:0] v1529; shift_adder #(7, 5, 1, 1, 8, 1, 1) op_1529 (v1403[6:0], v1373[4:0], v1529[7:0]); // 8.0
    wire [6:0] v1530; shift_adder #(5, 7, 1, 1, 7, -1, 0) op_1530 (v1405[4:0], v1392[6:0], v1530[6:0]); // 8.0
    wire [6:0] v1531; shift_adder #(5, 6, 0, 1, 7, 0, 1) op_1531 (v1406[4:0], v1407[5:0], v1531[6:0]); // 8.0
    wire [6:0] v1532; shift_adder #(6, 5, 1, 1, 7, 1, 0) op_1532 (v1408[5:0], v1409[4:0], v1532[6:0]); // 8.0
    wire [6:0] v1533; shift_adder #(5, 6, 1, 1, 7, 0, 0) op_1533 (v865[4:0], v1410[5:0], v1533[6:0]); // 8.0
    wire [7:0] v1534; shift_adder #(5, 7, 1, 1, 8, -1, 0) op_1534 (v1411[4:0], v1412[6:0], v1534[7:0]); // 8.0
    wire [7:0] v1535; shift_adder #(6, 5, 1, 1, 8, 2, 0) op_1535 (v1413[5:0], v1414[4:0], v1535[7:0]); // 8.0
    wire [7:0] v1536; shift_adder #(7, 6, 1, 1, 8, 0, 0) op_1536 (v1416[6:0], v1417[5:0], v1536[7:0]); // 8.0
    wire [6:0] v1537; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_1537 (v1418[5:0], v1419[5:0], v1537[6:0]); // 8.0
    wire [7:0] v1538; shift_adder #(7, 6, 1, 1, 8, 1, 0) op_1538 (v1267[6:0], v1420[5:0], v1538[7:0]); // 8.0
    wire [7:0] v1539; shift_adder #(7, 7, 1, 1, 8, 0, 0) op_1539 (v1421[6:0], v1422[6:0], v1539[7:0]); // 8.0
    wire [6:0] v1540; shift_adder #(5, 6, 1, 1, 7, 1, 1) op_1540 (v865[4:0], v1407[5:0], v1540[6:0]); // 8.0
    wire [6:0] v1541; shift_adder #(6, 5, 1, 1, 7, 0, 1) op_1541 (v1423[5:0], v1269[4:0], v1541[6:0]); // 8.0
    wire [6:0] v1542; shift_adder #(5, 6, 1, 1, 7, 0, 0) op_1542 (v1424[4:0], v1425[5:0], v1542[6:0]); // 8.0
    wire [6:0] v1543; shift_adder #(3, 6, 0, 1, 7, -2, 0) op_1543 (v1091[2:0], v1410[5:0], v1543[6:0]); // 8.0
    wire [6:0] v1544; shift_adder #(6, 6, 1, 1, 7, 0, 1) op_1544 (v1404[5:0], v1207[5:0], v1544[6:0]); // 8.0
    wire [6:0] v1545; shift_adder #(6, 7, 1, 1, 7, 0, 0) op_1545 (v1427[5:0], v1392[6:0], v1545[6:0]); // 8.0
    wire [5:0] v1546; shift_adder #(5, 4, 0, 1, 6, 0, 0) op_1546 (v1275[4:0], v1428[3:0], v1546[5:0]); // 8.0
    wire [7:0] v1547; shift_adder #(7, 5, 1, 1, 8, 2, 1) op_1547 (v1429[6:0], v1411[4:0], v1547[7:0]); // 8.0
    wire [7:0] v1548; shift_adder #(5, 7, 1, 1, 8, -1, 1) op_1548 (v1414[4:0], v1277[6:0], v1548[7:0]); // 8.0
    wire [6:0] v1549; shift_adder #(6, 4, 1, 1, 7, 1, 1) op_1549 (v1430[5:0], v1428[3:0], v1549[6:0]); // 8.0
    wire [5:0] v1550; shift_adder #(5, 6, 1, 1, 6, 0, 0) op_1550 (v1432[4:0], v1415[5:0], v1550[5:0]); // 8.0
    wire [6:0] v1551; shift_adder #(6, 6, 1, 1, 7, 0, 1) op_1551 (v1433[5:0], v1268[5:0], v1551[6:0]); // 8.0
    wire [7:0] v1552; shift_adder #(6, 5, 1, 0, 8, -1, 0) op_1552 (v1420[5:0], v1434[4:0], v1552[7:0]); // 8.0
    wire [7:0] v1553; shift_adder #(5, 7, 0, 1, 8, 0, 0) op_1553 (v1279[4:0], v1421[6:0], v1553[7:0]); // 8.0
    wire [5:0] v1554; shift_adder #(6, 5, 1, 1, 6, 0, 1) op_1554 (v1435[5:0], v1409[4:0], v1554[5:0]); // 8.0
    wire [7:0] v1555; shift_adder #(5, 7, 1, 1, 8, -1, 0) op_1555 (v1436[4:0], v1437[6:0], v1555[7:0]); // 8.0
    wire [6:0] v1556; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_1556 (v1438[4:0], v1439[4:0], v1556[6:0]); // 8.0
    wire [7:0] v1557; shift_adder #(7, 6, 1, 1, 8, 0, 0) op_1557 (v1441[6:0], v1442[5:0], v1557[7:0]); // 8.0
    wire [6:0] v1558; shift_adder #(6, 5, 1, 1, 7, 1, 0) op_1558 (v1443[5:0], v1444[4:0], v1558[6:0]); // 8.0
    wire [6:0] v1559; shift_adder #(7, 5, 1, 1, 7, 1, 1) op_1559 (v1445[6:0], v1446[4:0], v1559[6:0]); // 8.0
    wire [6:0] v1560; shift_adder #(5, 6, 1, 1, 7, 0, 1) op_1560 (v1439[4:0], v1298[5:0], v1560[6:0]); // 8.0
    wire [6:0] v1561; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_1561 (v1440[5:0], v1448[5:0], v1561[6:0]); // 8.0
    wire [6:0] v1562; shift_adder #(6, 5, 1, 1, 7, 0, 0) op_1562 (v1299[5:0], v1446[4:0], v1562[6:0]); // 8.0
    wire [6:0] v1563; shift_adder #(6, 5, 1, 1, 7, 1, 1) op_1563 (v1449[5:0], v1436[4:0], v1563[6:0]); // 8.0
    wire [7:0] v1564; shift_adder #(6, 7, 1, 1, 8, -1, 1) op_1564 (v1431[5:0], v1277[6:0], v1564[7:0]); // 8.0
    wire [6:0] v1565; shift_adder #(6, 6, 1, 1, 7, 1, 0) op_1565 (v1451[5:0], v1415[5:0], v1565[6:0]); // 8.0
    wire [5:0] v1566; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_1566 (v1452[4:0], v1453[4:0], v1566[5:0]); // 8.0
    wire [5:0] v1567; shift_adder #(4, 5, 0, 1, 6, 0, 0) op_1567 (v1307[3:0], v1454[4:0], v1567[5:0]); // 8.0
    wire [6:0] v1568; shift_adder #(7, 6, 1, 1, 7, 0, 1) op_1568 (v1455[6:0], v1456[5:0], v1568[6:0]); // 8.0
    wire [7:0] v1569; shift_adder #(4, 8, 1, 1, 8, -2, 0) op_1569 (v1457[3:0], v1458[7:0], v1569[7:0]); // 8.0
    wire [6:0] v1570; shift_adder #(5, 6, 1, 1, 7, 0, 1) op_1570 (v1452[4:0], v1317[5:0], v1570[6:0]); // 8.0
    wire [6:0] v1571; shift_adder #(6, 6, 1, 1, 7, 0, 1) op_1571 (v1447[5:0], v1298[5:0], v1571[6:0]); // 8.0
    wire [6:0] v1572; shift_adder #(6, 6, 1, 1, 7, 1, 0) op_1572 (v1461[5:0], v1440[5:0], v1572[6:0]); // 8.0
    wire [7:0] v1573; shift_adder #(7, 6, 1, 1, 8, 1, 0) op_1573 (v1462[6:0], v1463[5:0], v1573[7:0]); // 8.0
    wire [6:0] v1574; shift_adder #(6, 5, 1, 1, 7, 1, 0) op_1574 (v1464[5:0], v1453[4:0], v1574[6:0]); // 8.0
    wire [6:0] v1575; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_1575 (v1456[5:0], v1466[5:0], v1575[6:0]); // 8.0
    wire [6:0] v1576; shift_adder #(7, 4, 1, 1, 7, 2, 0) op_1576 (v1455[6:0], v1457[3:0], v1576[6:0]); // 8.0
    wire [7:0] v1577; shift_adder #(7, 6, 1, 1, 8, -1, 1) op_1577 (v1467[6:0], v1468[5:0], v1577[7:0]); // 8.0
    wire [4:0] v1578; shift_adder #(3, 5, 0, 1, 5, 0, 0) op_1578 (v937[2:0], v1469[4:0], v1578[4:0]); // 8.0
    wire [6:0] v1579; shift_adder #(4, 5, 0, 1, 7, -1, 0) op_1579 (v1307[3:0], v1470[4:0], v1579[6:0]); // 8.0
    wire [6:0] v1580; shift_adder #(6, 5, 1, 1, 7, 1, 1) op_1580 (v1471[5:0], v1148[4:0], v1580[6:0]); // 8.0
    wire [6:0] v1581; shift_adder #(6, 5, 0, 0, 7, 0, 0) op_1581 (v1472[5:0], v1473[4:0], v1581[6:0]); // 8.0
    wire [6:0] v1582; shift_adder #(4, 6, 0, 1, 7, -1, 0) op_1582 (v1332[3:0], v1471[5:0], v1582[6:0]); // 8.0
    wire [6:0] v1583; shift_adder #(4, 6, 0, 1, 7, -1, 0) op_1583 (v1475[3:0], v1476[5:0], v1583[6:0]); // 8.0
    wire [7:0] v1584; shift_adder #(5, 7, 1, 1, 8, -3, 0) op_1584 (v1333[4:0], v1478[6:0], v1584[7:0]); // 8.0
    wire [6:0] v1585; shift_adder #(6, 4, 0, 0, 7, 1, 1) op_1585 (v1479[5:0], v1332[3:0], v1585[6:0]); // 8.0
    wire [6:0] v1586; shift_adder #(6, 7, 1, 1, 7, -1, 1) op_1586 (v1480[5:0], v1467[6:0], v1586[6:0]); // 8.0
    wire [7:0] v1587; shift_adder #(6, 7, 1, 1, 8, 0, 1) op_1587 (v1468[5:0], v1339[6:0], v1587[7:0]); // 8.0
    wire [8:0] v1588; shift_adder #(6, 8, 1, 1, 9, -2, 0) op_1588 (v1340[5:0], v1482[7:0], v1588[8:0]); // 8.0
    wire [6:0] v1589; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_1589 (v1483[5:0], v1468[5:0], v1589[6:0]); // 8.0
    wire [6:0] v1590; shift_adder #(4, 5, 0, 1, 7, -1, 1) op_1590 (v1307[3:0], v1469[4:0], v1590[6:0]); // 8.0
    wire [5:0] v1591; shift_adder #(6, 5, 1, 1, 6, 1, 1) op_1591 (v1485[5:0], v1344[4:0], v1591[5:0]); // 8.0
    wire [7:0] v1592; shift_adder #(7, 8, 1, 1, 8, -1, 0) op_1592 (v1346[6:0], v1482[7:0], v1592[7:0]); // 8.0
    wire [7:0] v1593; shift_adder #(7, 6, 1, 1, 8, 1, 1) op_1593 (v1487[6:0], v1488[5:0], v1593[7:0]); // 8.0
    wire [7:0] v1594; shift_adder #(8, 2, 1, 0, 8, 0, 1) op_1594 (v1593[7:0], 2'b10, v1594[7:0]); // 8.0
    wire [6:0] v1595; assign v1595[6:0] = v1594[6:0] & {7{~v1594[7]}}; // 8.0
    wire [6:0] v1596; shift_adder #(7, 2, 0, 0, 7, 0, 0) op_1596 (v1595[6:0], 2'b10, v1596[6:0]); // 8.0
    wire [3:0] v1597; assign v1597[3:0] = v1596[5:2]; // 8.0
    wire [6:0] v1598; shift_adder #(6, 6, 1, 1, 7, 0, 0) op_1598 (v1490[5:0], v1491[5:0], v1598[6:0]); // 8.0
    wire [5:0] v1599; shift_adder #(5, 5, 1, 1, 6, -1, 0) op_1599 (v1353[4:0], v1493[4:0], v1599[5:0]); // 8.0
    wire [5:0] v1600; shift_adder #(6, 4, 1, 0, 6, 0, 1) op_1600 (v1495[5:0], v1351[3:0], v1600[5:0]); // 8.0
    wire [5:0] v1601; shift_adder #(5, 6, 1, 1, 6, 0, 1) op_1601 (v1496[4:0], v1488[5:0], v1601[5:0]); // 8.0
    wire [6:0] v1602; shift_adder #(7, 5, 1, 0, 7, 0, 1) op_1602 (v1497[6:0], v1357[4:0], v1602[6:0]); // 8.0
    wire [6:0] v1603; shift_adder #(6, 6, 1, 1, 7, 0, 1) op_1603 (v1465[5:0], v1317[5:0], v1603[6:0]); // 8.0
    wire [6:0] v1604; shift_adder #(6, 6, 1, 1, 7, 1, 0) op_1604 (v1499[5:0], v1456[5:0], v1604[6:0]); // 8.0
    wire [7:0] v1605; shift_adder #(6, 7, 1, 1, 8, -1, 0) op_1605 (v1362[5:0], v1501[6:0], v1605[7:0]); // 9.0
    wire [7:0] v1606; shift_adder #(7, 7, 1, 1, 8, 0, 0) op_1606 (v1502[6:0], v1503[6:0], v1606[7:0]); // 9.0
    wire [9:0] v1607; shift_adder #(8, 3, 1, 0, 10, -2, 1) op_1607 (v1606[7:0], 3'b101, v1607[9:0]); // 9.0
    wire [8:0] v1608; assign v1608[8:0] = v1607[8:0] & {9{~v1607[9]}}; // 9.0
    wire [8:0] v1609; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1609 (v1608[8:0], 3'b100, v1609[8:0]); // 9.0
    wire [4:0] v1610; assign v1610[4:0] = v1609[7:3]; // 9.0
    wire [6:0] v1611; shift_adder #(7, 5, 1, 1, 7, 0, 1) op_1611 (v1505[6:0], v1372[4:0], v1611[6:0]); // 9.0
    wire [7:0] v1612; shift_adder #(7, 7, 1, 1, 8, 0, 0) op_1612 (v1507[6:0], v1508[6:0], v1612[7:0]); // 9.0
    wire [6:0] v1613; shift_adder #(7, 6, 1, 1, 7, 0, 0) op_1613 (v1509[6:0], v1510[5:0], v1613[6:0]); // 9.0
    wire [7:0] v1614; shift_adder #(7, 7, 1, 1, 8, 0, 0) op_1614 (v1513[6:0], v1514[6:0], v1614[7:0]); // 9.0
    wire [7:0] v1615; shift_adder #(8, 6, 1, 1, 8, 1, 1) op_1615 (v1516[7:0], v1386[5:0], v1615[7:0]); // 9.0
    wire [7:0] v1616; shift_adder #(8, 7, 1, 1, 8, 0, 0) op_1616 (v1388[7:0], v1518[6:0], v1616[7:0]); // 9.0
    wire [7:0] v1617; shift_adder #(7, 7, 1, 1, 8, -1, 1) op_1617 (v1520[6:0], v1392[6:0], v1617[7:0]); // 9.0
    wire [6:0] v1618; shift_adder #(7, 5, 1, 1, 7, 0, 1) op_1618 (v1522[6:0], v1376[4:0], v1618[6:0]); // 9.0
    wire [7:0] v1619; shift_adder #(7, 6, 1, 1, 8, 1, 1) op_1619 (v1523[6:0], v1387[5:0], v1619[7:0]); // 9.0
    wire [7:0] v1620; shift_adder #(6, 7, 1, 1, 8, 0, 0) op_1620 (v1524[5:0], v1514[6:0], v1620[7:0]); // 9.0
    wire [8:0] v1621; shift_adder #(7, 8, 1, 1, 9, 0, 0) op_1621 (v1525[6:0], v1526[7:0], v1621[8:0]); // 9.0
    wire [8:0] v1622; shift_adder #(9, 2, 1, 0, 9, 0, 1) op_1622 (v1621[8:0], 2'b10, v1622[8:0]); // 9.0
    wire [7:0] v1623; assign v1623[7:0] = v1622[7:0] & {8{~v1622[8]}}; // 9.0
    wire [7:0] v1624; shift_adder #(8, 2, 0, 0, 8, 0, 0) op_1624 (v1623[7:0], 2'b10, v1624[7:0]); // 9.0
    wire [3:0] v1625; assign v1625[3:0] = v1624[5:2]; // 9.0
    wire [7:0] v1626; shift_adder #(7, 7, 1, 1, 8, 0, 0) op_1626 (v1527[6:0], v1528[6:0], v1626[7:0]); // 9.0
    wire [7:0] v1627; shift_adder #(8, 2, 1, 0, 8, 0, 0) op_1627 (v1626[7:0], 2'b10, v1627[7:0]); // 9.0
    wire [6:0] v1628; assign v1628[6:0] = v1627[6:0] & {7{~v1627[7]}}; // 9.0
    wire [6:0] v1629; shift_adder #(7, 2, 0, 0, 7, 0, 0) op_1629 (v1628[6:0], 2'b10, v1629[6:0]); // 9.0
    wire [3:0] v1630; assign v1630[3:0] = v1629[5:2]; // 9.0
    wire [8:0] v1631; shift_adder #(8, 6, 1, 1, 9, 2, 1) op_1631 (v1529[7:0], v1404[5:0], v1631[8:0]); // 9.0
    wire [8:0] v1632; shift_adder #(7, 7, 1, 1, 9, 1, 0) op_1632 (v1530[6:0], v1508[6:0], v1632[8:0]); // 9.0
    wire [7:0] v1633; shift_adder #(7, 7, 1, 1, 8, 0, 0) op_1633 (v1532[6:0], v1533[6:0], v1633[7:0]); // 9.0
    wire [7:0] v1634; shift_adder #(8, 6, 1, 1, 8, 1, 1) op_1634 (v1535[7:0], v1415[5:0], v1634[7:0]); // 9.0
    wire [6:0] v1635; shift_adder #(7, 5, 1, 1, 7, 0, 1) op_1635 (v1537[6:0], v1414[4:0], v1635[6:0]); // 9.0
    wire [8:0] v1636; shift_adder #(8, 8, 1, 1, 9, 1, 0) op_1636 (v1538[7:0], v1539[7:0], v1636[8:0]); // 9.0
    wire [7:0] v1637; shift_adder #(7, 7, 1, 1, 8, 1, 0) op_1637 (v1541[6:0], v1542[6:0], v1637[7:0]); // 9.0
    wire [7:0] v1638; shift_adder #(8, 7, 1, 1, 8, 0, 0) op_1638 (v1426[7:0], v1545[6:0], v1638[7:0]); // 9.0
    wire [8:0] v1639; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_1639 (v1547[7:0], v1548[7:0], v1639[8:0]); // 9.0
    wire [7:0] v1640; shift_adder #(7, 6, 1, 1, 8, 1, 1) op_1640 (v1549[6:0], v1431[5:0], v1640[7:0]); // 9.0
    wire [8:0] v1641; shift_adder #(6, 8, 1, 1, 9, -1, 0) op_1641 (v1550[5:0], v1548[7:0], v1641[8:0]); // 9.0
    wire [7:0] v1642; shift_adder #(7, 7, 1, 1, 8, 1, 0) op_1642 (v1543[6:0], v1551[6:0], v1642[7:0]); // 9.0
    wire [8:0] v1643; shift_adder #(8, 7, 1, 1, 9, -1, 0) op_1643 (v1552[7:0], v1540[6:0], v1643[8:0]); // 9.0
    wire [8:0] v1644; shift_adder #(7, 6, 1, 1, 9, 2, 0) op_1644 (v1533[6:0], v1554[5:0], v1644[8:0]); // 9.0
    wire [6:0] v1645; shift_adder #(7, 6, 1, 1, 7, 0, 1) op_1645 (v1556[6:0], v1440[5:0], v1645[6:0]); // 9.0
    wire [6:0] v1646; shift_adder #(7, 5, 1, 1, 7, 0, 1) op_1646 (v1558[6:0], v1439[4:0], v1646[6:0]); // 9.0
    wire [8:0] v1647; shift_adder #(7, 6, 1, 1, 9, 2, 1) op_1647 (v1559[6:0], v1447[5:0], v1647[8:0]); // 9.0
    wire [7:0] v1648; shift_adder #(7, 7, 1, 1, 8, 0, 0) op_1648 (v1560[6:0], v1561[6:0], v1648[7:0]); // 9.0
    wire [7:0] v1649; shift_adder #(7, 7, 1, 1, 8, 0, 0) op_1649 (v1563[6:0], v1560[6:0], v1649[7:0]); // 9.0
    wire [8:0] v1650; shift_adder #(8, 7, 1, 1, 9, 0, 0) op_1650 (v1450[7:0], v1565[6:0], v1650[8:0]); // 9.0
    wire [7:0] v1651; shift_adder #(6, 7, 1, 1, 8, 0, 0) op_1651 (v1567[5:0], v1568[6:0], v1651[7:0]); // 9.0
    wire [7:0] v1652; shift_adder #(7, 7, 1, 1, 8, 0, 1) op_1652 (v1570[6:0], v1459[6:0], v1652[7:0]); // 9.0
    wire [7:0] v1653; shift_adder #(8, 7, 1, 1, 8, 0, 0) op_1653 (v1460[7:0], v1572[6:0], v1653[7:0]); // 9.0
    wire [6:0] v1654; shift_adder #(7, 5, 1, 1, 7, 0, 1) op_1654 (v1574[6:0], v1452[4:0], v1654[6:0]); // 9.0
    wire [7:0] v1655; shift_adder #(7, 6, 1, 1, 8, 1, 1) op_1655 (v1570[6:0], v1465[5:0], v1655[7:0]); // 9.0
    wire [7:0] v1656; shift_adder #(7, 7, 1, 1, 8, -1, 1) op_1656 (v1575[6:0], v1576[6:0], v1656[7:0]); // 9.0
    wire [6:0] v1657; shift_adder #(5, 7, 1, 1, 7, -1, 0) op_1657 (v1578[4:0], v1579[6:0], v1657[6:0]); // 9.0
    wire [8:0] v1658; shift_adder #(7, 7, 1, 0, 9, 1, 1) op_1658 (v1580[6:0], v1581[6:0], v1658[8:0]); // 9.0
    wire [9:0] v1659; shift_adder #(9, 4, 1, 0, 10, -1, 0) op_1659 (v1658[8:0], 4'b1011, v1659[9:0]); // 9.0
    wire [6:0] v1660; assign v1660[6:0] = v1659[6:0] & {7{~v1659[9]}}; // 9.0
    wire [6:0] v1661; shift_adder #(7, 4, 0, 0, 7, 0, 0) op_1661 (v1660[6:0], 4'b1000, v1661[6:0]); // 9.0
    wire [2:0] v1662; assign v1662[2:0] = v1661[6:4]; // 9.0
    wire [7:0] v1663; shift_adder #(7, 7, 1, 1, 8, 0, 0) op_1663 (v1474[6:0], v1582[6:0], v1663[7:0]); // 9.0
    wire [9:0] v1664; shift_adder #(8, 4, 1, 0, 10, -2, 1) op_1664 (v1663[7:0], 4'b1001, v1664[9:0]); // 9.0
    wire [8:0] v1665; assign v1665[8:0] = v1664[8:0] & {9{~v1664[9]}}; // 9.0
    wire [8:0] v1666; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1666 (v1665[8:0], 3'b100, v1666[8:0]); // 9.0
    wire [4:0] v1667; assign v1667[4:0] = v1666[7:3]; // 9.0
    wire [7:0] v1668; shift_adder #(7, 6, 1, 1, 8, -1, 1) op_1668 (v1583[6:0], v1471[5:0], v1668[7:0]); // 9.0
    wire [8:0] v1669; shift_adder #(8, 3, 1, 0, 9, -1, 1) op_1669 (v1668[7:0], 3'b101, v1669[8:0]); // 9.0
    wire [7:0] v1670; assign v1670[7:0] = v1669[7:0] & {8{~v1669[8]}}; // 9.0
    wire [7:0] v1671; shift_adder #(8, 3, 0, 0, 8, 0, 0) op_1671 (v1670[7:0], 3'b100, v1671[7:0]); // 9.0
    wire [4:0] v1672; assign v1672[4:0] = v1671[7:3]; // 9.0
    wire [8:0] v1673; shift_adder #(7, 8, 1, 1, 9, -1, 0) op_1673 (v1477[6:0], v1584[7:0], v1673[8:0]); // 9.0
    wire [8:0] v1674; shift_adder #(9, 3, 1, 0, 9, 0, 1) op_1674 (v1673[8:0], 3'b100, v1674[8:0]); // 9.0
    wire [7:0] v1675; assign v1675[7:0] = v1674[7:0] & {8{~v1674[8]}}; // 9.0
    wire [7:0] v1676; shift_adder #(8, 2, 0, 0, 8, 0, 0) op_1676 (v1675[7:0], 2'b10, v1676[7:0]); // 9.0
    wire [4:0] v1677; assign v1677[4:0] = v1676[6:2]; // 9.0
    wire [7:0] v1678; shift_adder #(7, 7, 1, 1, 8, 1, 0) op_1678 (v1580[6:0], v1585[6:0], v1678[7:0]); // 9.0
    wire [8:0] v1679; shift_adder #(8, 3, 1, 0, 9, 0, 0) op_1679 (v1678[7:0], 3'b100, v1679[8:0]); // 9.0
    wire [7:0] v1680; assign v1680[7:0] = v1679[7:0] & {8{~v1679[8]}}; // 9.0
    wire [7:0] v1681; shift_adder #(8, 2, 0, 0, 8, 0, 0) op_1681 (v1680[7:0], 2'b10, v1681[7:0]); // 9.0
    wire [4:0] v1682; assign v1682[4:0] = v1681[6:2]; // 9.0
    wire [8:0] v1683; shift_adder #(7, 8, 1, 1, 9, 0, 0) op_1683 (v1586[6:0], v1587[7:0], v1683[8:0]); // 9.0
    wire [6:0] v1684; shift_adder #(5, 5, 1, 0, 7, 1, 1) op_1684 (v1578[4:0], v1481[4:0], v1684[6:0]); // 9.0
    wire [7:0] v1685; shift_adder #(5, 7, 0, 1, 8, 0, 0) op_1685 (v1481[4:0], v1589[6:0], v1685[7:0]); // 9.0
    wire [8:0] v1686; shift_adder #(8, 6, 1, 1, 9, 1, 0) op_1686 (v1484[7:0], v1591[5:0], v1686[8:0]); // 9.0
    wire [8:0] v1687; shift_adder #(6, 8, 1, 1, 9, -1, 0) op_1687 (v1486[5:0], v1592[7:0], v1687[8:0]); // 9.0
    wire [7:0] v1688; shift_adder #(5, 7, 0, 1, 8, 0, 0) op_1688 (v1489[4:0], v1598[6:0], v1688[7:0]); // 9.0
    wire [9:0] v1689; shift_adder #(8, 4, 1, 0, 10, -2, 1) op_1689 (v1688[7:0], 4'b1001, v1689[9:0]); // 9.0
    wire [8:0] v1690; assign v1690[8:0] = v1689[8:0] & {9{~v1689[9]}}; // 9.0
    wire [8:0] v1691; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1691 (v1690[8:0], 3'b100, v1691[8:0]); // 9.0
    wire [4:0] v1692; assign v1692[4:0] = v1691[7:3]; // 9.0
    wire [7:0] v1693; shift_adder #(7, 6, 1, 1, 8, 0, 0) op_1693 (v1492[6:0], v1599[5:0], v1693[7:0]); // 9.0
    wire [9:0] v1694; shift_adder #(8, 3, 1, 0, 10, -2, 1) op_1694 (v1693[7:0], 3'b101, v1694[9:0]); // 9.0
    wire [8:0] v1695; assign v1695[8:0] = v1694[8:0] & {9{~v1694[9]}}; // 9.0
    wire [8:0] v1696; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1696 (v1695[8:0], 3'b100, v1696[8:0]); // 9.0
    wire [4:0] v1697; assign v1697[4:0] = v1696[7:3]; // 9.0
    wire [6:0] v1698; shift_adder #(7, 6, 1, 1, 7, 1, 0) op_1698 (v1494[6:0], v1600[5:0], v1698[6:0]); // 9.0
    wire [6:0] v1699; shift_adder #(7, 2, 1, 0, 7, 0, 0) op_1699 (v1698[6:0], 2'b10, v1699[6:0]); // 9.0
    wire [5:0] v1700; assign v1700[5:0] = v1699[5:0] & {6{~v1699[6]}}; // 9.0
    wire [5:0] v1701; shift_adder #(6, 2, 0, 0, 6, 0, 0) op_1701 (v1700[5:0], 2'b10, v1701[5:0]); // 9.0
    wire [3:0] v1702; assign v1702[3:0] = v1701[5:2]; // 9.0
    wire [7:0] v1703; shift_adder #(6, 7, 1, 1, 8, 0, 0) op_1703 (v1601[5:0], v1602[6:0], v1703[7:0]); // 9.0
    wire [9:0] v1704; shift_adder #(8, 4, 1, 0, 10, -2, 0) op_1704 (v1703[7:0], 4'b1011, v1704[9:0]); // 9.0
    wire [7:0] v1705; assign v1705[7:0] = v1704[7:0] & {8{~v1704[9]}}; // 9.0
    wire [7:0] v1706; shift_adder #(8, 3, 0, 0, 8, 0, 0) op_1706 (v1705[7:0], 3'b100, v1706[7:0]); // 9.0
    wire [4:0] v1707; assign v1707[4:0] = v1706[7:3]; // 9.0
    wire [7:0] v1708; shift_adder #(8, 7, 1, 1, 8, 0, 0) op_1708 (v1498[7:0], v1604[6:0], v1708[7:0]); // 9.0
    wire [8:0] v1709; shift_adder #(8, 8, 1, 1, 9, 1, 0) op_1709 (v1500[7:0], v1605[7:0], v1709[8:0]); // 10.0
    wire [9:0] v1710; shift_adder #(9, 4, 1, 0, 10, -1, 1) op_1710 (v1709[8:0], 4'b1001, v1710[9:0]); // 10.0
    wire [8:0] v1711; assign v1711[8:0] = v1710[8:0] & {9{~v1710[9]}}; // 10.0
    wire [8:0] v1712; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1712 (v1711[8:0], 3'b100, v1712[8:0]); // 10.0
    wire [4:0] v1713; assign v1713[4:0] = v1712[7:3]; // 10.0
    wire [8:0] v1714; shift_adder #(8, 7, 1, 1, 9, 0, 0) op_1714 (v1504[7:0], v1611[6:0], v1714[8:0]); // 10.0
    wire [9:0] v1715; shift_adder #(9, 3, 1, 0, 10, -2, 1) op_1715 (v1714[8:0], 3'b101, v1715[9:0]); // 10.0
    wire [8:0] v1716; assign v1716[8:0] = v1715[8:0] & {9{~v1715[9]}}; // 10.0
    wire [8:0] v1717; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1717 (v1716[8:0], 3'b100, v1717[8:0]); // 10.0
    wire [5:0] v1718; assign v1718[5:0] = v1717[8:3]; // 10.0
    wire [7:0] v1719; shift_adder #(7, 8, 1, 1, 8, 0, 0) op_1719 (v1506[6:0], v1612[7:0], v1719[7:0]); // 10.0
    wire [7:0] v1720; shift_adder #(8, 2, 1, 0, 8, 0, 0) op_1720 (v1719[7:0], 2'b10, v1720[7:0]); // 10.0
    wire [6:0] v1721; assign v1721[6:0] = v1720[6:0] & {7{~v1720[7]}}; // 10.0
    wire [6:0] v1722; shift_adder #(7, 1, 0, 0, 7, 0, 0) op_1722 (v1721[6:0], 1'b1, v1722[6:0]); // 10.0
    wire [4:0] v1723; assign v1723[4:0] = v1722[5:1]; // 10.0
    wire [7:0] v1724; shift_adder #(7, 8, 1, 1, 8, 0, 1) op_1724 (v1613[6:0], v1511[7:0], v1724[7:0]); // 10.0
    wire [9:0] v1725; shift_adder #(8, 4, 1, 0, 10, -2, 0) op_1725 (v1724[7:0], 4'b1011, v1725[9:0]); // 10.0
    wire [8:0] v1726; assign v1726[8:0] = v1725[8:0] & {9{~v1725[9]}}; // 10.0
    wire [8:0] v1727; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1727 (v1726[8:0], 3'b100, v1727[8:0]); // 10.0
    wire [4:0] v1728; assign v1728[4:0] = v1727[7:3]; // 10.0
    wire [7:0] v1729; shift_adder #(7, 8, 1, 1, 8, 0, 0) op_1729 (v1512[6:0], v1614[7:0], v1729[7:0]); // 10.0
    wire [7:0] v1730; shift_adder #(8, 2, 1, 0, 8, 0, 0) op_1730 (v1729[7:0], 2'b10, v1730[7:0]); // 10.0
    wire [6:0] v1731; assign v1731[6:0] = v1730[6:0] & {7{~v1730[7]}}; // 10.0
    wire [6:0] v1732; shift_adder #(7, 2, 0, 0, 7, 0, 0) op_1732 (v1731[6:0], 2'b10, v1732[6:0]); // 10.0
    wire [3:0] v1733; assign v1733[3:0] = v1732[5:2]; // 10.0
    wire [8:0] v1734; shift_adder #(8, 8, 1, 1, 9, -1, 0) op_1734 (v1515[7:0], v1615[7:0], v1734[8:0]); // 10.0
    wire [9:0] v1735; shift_adder #(9, 4, 1, 0, 10, -1, 1) op_1735 (v1734[8:0], 4'b1001, v1735[9:0]); // 10.0
    wire [8:0] v1736; assign v1736[8:0] = v1735[8:0] & {9{~v1735[9]}}; // 10.0
    wire [8:0] v1737; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1737 (v1736[8:0], 3'b100, v1737[8:0]); // 10.0
    wire [4:0] v1738; assign v1738[4:0] = v1737[7:3]; // 10.0
    wire [8:0] v1739; shift_adder #(7, 8, 1, 1, 9, 0, 0) op_1739 (v1517[6:0], v1616[7:0], v1739[8:0]); // 10.0
    wire [8:0] v1740; shift_adder #(9, 2, 1, 0, 9, 0, 1) op_1740 (v1739[8:0], 2'b10, v1740[8:0]); // 10.0
    wire [7:0] v1741; assign v1741[7:0] = v1740[7:0] & {8{~v1740[8]}}; // 10.0
    wire [7:0] v1742; shift_adder #(8, 1, 0, 0, 8, 0, 0) op_1742 (v1741[7:0], 1'b1, v1742[7:0]); // 10.0
    wire [4:0] v1743; assign v1743[4:0] = v1742[5:1]; // 10.0
    wire [8:0] v1744; shift_adder #(8, 8, 1, 1, 9, -1, 0) op_1744 (v1519[7:0], v1617[7:0], v1744[8:0]); // 10.0
    wire [9:0] v1745; shift_adder #(9, 4, 1, 0, 10, -1, 1) op_1745 (v1744[8:0], 4'b1001, v1745[9:0]); // 10.0
    wire [8:0] v1746; assign v1746[8:0] = v1745[8:0] & {9{~v1745[9]}}; // 10.0
    wire [8:0] v1747; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1747 (v1746[8:0], 3'b100, v1747[8:0]); // 10.0
    wire [4:0] v1748; assign v1748[4:0] = v1747[7:3]; // 10.0
    wire [9:0] v1749; shift_adder #(9, 7, 1, 1, 10, 1, 0) op_1749 (v1521[8:0], v1618[6:0], v1749[9:0]); // 10.0
    wire [9:0] v1750; shift_adder #(10, 3, 1, 0, 10, -1, 1) op_1750 (v1749[9:0], 3'b101, v1750[9:0]); // 10.0
    wire [8:0] v1751; assign v1751[8:0] = v1750[8:0] & {9{~v1750[9]}}; // 10.0
    wire [9:0] v1752; shift_adder #(9, 3, 0, 0, 10, 0, 0) op_1752 (v1751[8:0], 3'b100, v1752[9:0]); // 10.0
    wire [4:0] v1753; assign v1753[4:0] = v1752[7:3]; // 10.0
    wire [8:0] v1754; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_1754 (v1619[7:0], v1620[7:0], v1754[8:0]); // 10.0
    wire [10:0] v1755; shift_adder #(9, 4, 1, 0, 11, -2, 0) op_1755 (v1754[8:0], 4'b1011, v1755[10:0]); // 10.0
    wire [8:0] v1756; assign v1756[8:0] = v1755[8:0] & {9{~v1755[10]}}; // 10.0
    wire [8:0] v1757; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1757 (v1756[8:0], 3'b100, v1757[8:0]); // 10.0
    wire [4:0] v1758; assign v1758[4:0] = v1757[7:3]; // 10.0
    wire [5:0] v1759; shift_adder #(4, 4, 1, 1, 6, -1, 0) op_1759 (v1625[3:0], v1630[3:0], v1759[5:0]); // 10.0
    wire [9:0] v1760; shift_adder #(9, 9, 1, 1, 10, 0, 0) op_1760 (v1631[8:0], v1632[8:0], v1760[9:0]); // 10.0
    wire [10:0] v1761; shift_adder #(10, 4, 1, 0, 11, -1, 0) op_1761 (v1760[9:0], 4'b1011, v1761[10:0]); // 10.0
    wire [8:0] v1762; assign v1762[8:0] = v1761[8:0] & {9{~v1761[10]}}; // 10.0
    wire [8:0] v1763; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1763 (v1762[8:0], 3'b100, v1763[8:0]); // 10.0
    wire [4:0] v1764; assign v1764[4:0] = v1763[7:3]; // 10.0
    wire [7:0] v1765; shift_adder #(7, 8, 1, 1, 8, 0, 0) op_1765 (v1531[6:0], v1633[7:0], v1765[7:0]); // 10.0
    wire [9:0] v1766; shift_adder #(8, 4, 1, 0, 10, -2, 1) op_1766 (v1765[7:0], 4'b1001, v1766[9:0]); // 10.0
    wire [8:0] v1767; assign v1767[8:0] = v1766[8:0] & {9{~v1766[9]}}; // 10.0
    wire [8:0] v1768; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1768 (v1767[8:0], 3'b100, v1768[8:0]); // 10.0
    wire [4:0] v1769; assign v1769[4:0] = v1768[7:3]; // 10.0
    wire [8:0] v1770; shift_adder #(8, 8, 1, 1, 9, -1, 0) op_1770 (v1534[7:0], v1634[7:0], v1770[8:0]); // 10.0
    wire [9:0] v1771; shift_adder #(9, 4, 1, 0, 10, -1, 1) op_1771 (v1770[8:0], 4'b1001, v1771[9:0]); // 10.0
    wire [8:0] v1772; assign v1772[8:0] = v1771[8:0] & {9{~v1771[9]}}; // 10.0
    wire [8:0] v1773; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1773 (v1772[8:0], 3'b100, v1773[8:0]); // 10.0
    wire [5:0] v1774; assign v1774[5:0] = v1773[8:3]; // 10.0
    wire [8:0] v1775; shift_adder #(8, 7, 1, 1, 9, 0, 0) op_1775 (v1536[7:0], v1635[6:0], v1775[8:0]); // 10.0
    wire [9:0] v1776; shift_adder #(9, 3, 1, 0, 10, -2, 1) op_1776 (v1775[8:0], 3'b101, v1776[9:0]); // 10.0
    wire [8:0] v1777; assign v1777[8:0] = v1776[8:0] & {9{~v1776[9]}}; // 10.0
    wire [9:0] v1778; shift_adder #(9, 3, 0, 0, 10, 0, 0) op_1778 (v1777[8:0], 3'b100, v1778[9:0]); // 10.0
    wire [5:0] v1779; assign v1779[5:0] = v1778[8:3]; // 10.0
    wire [9:0] v1780; shift_adder #(9, 7, 1, 1, 10, 1, 1) op_1780 (v1636[8:0], v1540[6:0], v1780[9:0]); // 10.0
    wire [9:0] v1781; shift_adder #(10, 3, 1, 0, 10, 0, 1) op_1781 (v1780[9:0], 3'b100, v1781[9:0]); // 10.0
    wire [8:0] v1782; assign v1782[8:0] = v1781[8:0] & {9{~v1781[9]}}; // 10.0
    wire [8:0] v1783; shift_adder #(9, 2, 0, 0, 9, 0, 0) op_1783 (v1782[8:0], 2'b10, v1783[8:0]); // 10.0
    wire [4:0] v1784; assign v1784[4:0] = v1783[6:2]; // 10.0
    wire [9:0] v1785; shift_adder #(8, 7, 1, 1, 10, -1, 1) op_1785 (v1637[7:0], v1543[6:0], v1785[9:0]); // 10.0
    wire [9:0] v1786; shift_adder #(10, 3, 1, 0, 10, -1, 1) op_1786 (v1785[9:0], 3'b101, v1786[9:0]); // 10.0
    wire [8:0] v1787; assign v1787[8:0] = v1786[8:0] & {9{~v1786[9]}}; // 10.0
    wire [8:0] v1788; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1788 (v1787[8:0], 3'b100, v1788[8:0]); // 10.0
    wire [5:0] v1789; assign v1789[5:0] = v1788[8:3]; // 10.0
    wire [8:0] v1790; shift_adder #(7, 8, 1, 1, 9, 0, 0) op_1790 (v1544[6:0], v1638[7:0], v1790[8:0]); // 10.0
    wire [8:0] v1791; shift_adder #(9, 2, 1, 0, 9, 0, 1) op_1791 (v1790[8:0], 2'b10, v1791[8:0]); // 10.0
    wire [7:0] v1792; assign v1792[7:0] = v1791[7:0] & {8{~v1791[8]}}; // 10.0
    wire [7:0] v1793; shift_adder #(8, 1, 0, 0, 8, 0, 0) op_1793 (v1792[7:0], 1'b1, v1793[7:0]); // 10.0
    wire [5:0] v1794; assign v1794[5:0] = v1793[6:1]; // 10.0
    wire [8:0] v1795; shift_adder #(6, 9, 1, 1, 9, -2, 0) op_1795 (v1546[5:0], v1639[8:0], v1795[8:0]); // 10.0
    wire [8:0] v1796; shift_adder #(9, 3, 1, 0, 9, 0, 0) op_1796 (v1795[8:0], 3'b100, v1796[8:0]); // 10.0
    wire [7:0] v1797; assign v1797[7:0] = v1796[7:0] & {8{~v1796[8]}}; // 10.0
    wire [7:0] v1798; shift_adder #(8, 2, 0, 0, 8, 0, 0) op_1798 (v1797[7:0], 2'b10, v1798[7:0]); // 10.0
    wire [4:0] v1799; assign v1799[4:0] = v1798[6:2]; // 10.0
    wire [9:0] v1800; shift_adder #(8, 9, 1, 1, 10, -1, 0) op_1800 (v1640[7:0], v1641[8:0], v1800[9:0]); // 10.0
    wire [10:0] v1801; shift_adder #(10, 4, 1, 0, 11, -1, 0) op_1801 (v1800[9:0], 4'b1011, v1801[10:0]); // 10.0
    wire [8:0] v1802; assign v1802[8:0] = v1801[8:0] & {9{~v1801[10]}}; // 10.0
    wire [8:0] v1803; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1803 (v1802[8:0], 3'b100, v1803[8:0]); // 10.0
    wire [4:0] v1804; assign v1804[4:0] = v1803[7:3]; // 10.0
    wire [9:0] v1805; shift_adder #(8, 9, 1, 1, 10, 0, 1) op_1805 (v1642[7:0], v1643[8:0], v1805[9:0]); // 10.0
    wire [10:0] v1806; shift_adder #(10, 4, 1, 0, 11, -1, 0) op_1806 (v1805[9:0], 4'b1011, v1806[10:0]); // 10.0
    wire [8:0] v1807; assign v1807[8:0] = v1806[8:0] & {9{~v1806[10]}}; // 10.0
    wire [8:0] v1808; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1808 (v1807[8:0], 3'b100, v1808[8:0]); // 10.0
    wire [4:0] v1809; assign v1809[4:0] = v1808[7:3]; // 10.0
    wire [8:0] v1810; shift_adder #(8, 9, 1, 1, 9, -1, 0) op_1810 (v1553[7:0], v1644[8:0], v1810[8:0]); // 10.0
    wire [8:0] v1811; shift_adder #(9, 3, 1, 0, 9, 0, 0) op_1811 (v1810[8:0], 3'b100, v1811[8:0]); // 10.0
    wire [7:0] v1812; assign v1812[7:0] = v1811[7:0] & {8{~v1811[8]}}; // 10.0
    wire [7:0] v1813; shift_adder #(8, 2, 0, 0, 8, 0, 0) op_1813 (v1812[7:0], 2'b10, v1813[7:0]); // 10.0
    wire [4:0] v1814; assign v1814[4:0] = v1813[6:2]; // 10.0
    wire [7:0] v1815; shift_adder #(8, 7, 1, 1, 8, 0, 0) op_1815 (v1555[7:0], v1645[6:0], v1815[7:0]); // 10.0
    wire [9:0] v1816; shift_adder #(8, 4, 1, 0, 10, -2, 1) op_1816 (v1815[7:0], 4'b1001, v1816[9:0]); // 10.0
    wire [8:0] v1817; assign v1817[8:0] = v1816[8:0] & {9{~v1816[9]}}; // 10.0
    wire [8:0] v1818; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1818 (v1817[8:0], 3'b100, v1818[8:0]); // 10.0
    wire [5:0] v1819; assign v1819[5:0] = v1818[8:3]; // 10.0
    wire [7:0] v1820; shift_adder #(8, 7, 1, 1, 8, 0, 0) op_1820 (v1557[7:0], v1646[6:0], v1820[7:0]); // 10.0
    wire [9:0] v1821; shift_adder #(8, 3, 1, 0, 10, -2, 1) op_1821 (v1820[7:0], 3'b101, v1821[9:0]); // 10.0
    wire [8:0] v1822; assign v1822[8:0] = v1821[8:0] & {9{~v1821[9]}}; // 10.0
    wire [8:0] v1823; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1823 (v1822[8:0], 3'b100, v1823[8:0]); // 10.0
    wire [5:0] v1824; assign v1824[5:0] = v1823[8:3]; // 10.0
    wire [9:0] v1825; shift_adder #(9, 8, 1, 1, 10, 1, 0) op_1825 (v1647[8:0], v1648[7:0], v1825[9:0]); // 10.0
    wire [10:0] v1826; shift_adder #(10, 4, 1, 0, 11, -1, 0) op_1826 (v1825[9:0], 4'b1011, v1826[10:0]); // 10.0
    wire [8:0] v1827; assign v1827[8:0] = v1826[8:0] & {9{~v1826[10]}}; // 10.0
    wire [8:0] v1828; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1828 (v1827[8:0], 3'b100, v1828[8:0]); // 10.0
    wire [4:0] v1829; assign v1829[4:0] = v1828[7:3]; // 10.0
    wire [7:0] v1830; shift_adder #(7, 8, 1, 1, 8, 0, 0) op_1830 (v1562[6:0], v1649[7:0], v1830[7:0]); // 10.0
    wire [7:0] v1831; shift_adder #(8, 2, 1, 0, 8, 0, 0) op_1831 (v1830[7:0], 2'b10, v1831[7:0]); // 10.0
    wire [6:0] v1832; assign v1832[6:0] = v1831[6:0] & {7{~v1831[7]}}; // 10.0
    wire [6:0] v1833; shift_adder #(7, 1, 0, 0, 7, 0, 0) op_1833 (v1832[6:0], 1'b1, v1833[6:0]); // 10.0
    wire [4:0] v1834; assign v1834[4:0] = v1833[5:1]; // 10.0
    wire [9:0] v1835; shift_adder #(8, 9, 1, 1, 10, 1, 0) op_1835 (v1564[7:0], v1650[8:0], v1835[9:0]); // 10.0
    wire [9:0] v1836; shift_adder #(10, 3, 1, 0, 10, 0, 1) op_1836 (v1835[9:0], 3'b100, v1836[9:0]); // 10.0
    wire [8:0] v1837; assign v1837[8:0] = v1836[8:0] & {9{~v1836[9]}}; // 10.0
    wire [8:0] v1838; shift_adder #(9, 2, 0, 0, 9, 0, 0) op_1838 (v1837[8:0], 2'b10, v1838[8:0]); // 10.0
    wire [4:0] v1839; assign v1839[4:0] = v1838[6:2]; // 10.0
    wire [7:0] v1840; shift_adder #(6, 8, 1, 1, 8, -1, 0) op_1840 (v1566[5:0], v1651[7:0], v1840[7:0]); // 10.0
    wire [9:0] v1841; shift_adder #(8, 4, 1, 0, 10, -2, 1) op_1841 (v1840[7:0], 4'b1001, v1841[9:0]); // 10.0
    wire [8:0] v1842; assign v1842[8:0] = v1841[8:0] & {9{~v1841[9]}}; // 10.0
    wire [8:0] v1843; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1843 (v1842[8:0], 3'b100, v1843[8:0]); // 10.0
    wire [4:0] v1844; assign v1844[4:0] = v1843[7:3]; // 10.0
    wire [8:0] v1845; shift_adder #(8, 8, 1, 1, 9, 1, 0) op_1845 (v1569[7:0], v1652[7:0], v1845[8:0]); // 10.0
    wire [8:0] v1846; shift_adder #(9, 3, 1, 0, 9, 0, 0) op_1846 (v1845[8:0], 3'b100, v1846[8:0]); // 10.0
    wire [7:0] v1847; assign v1847[7:0] = v1846[7:0] & {8{~v1846[8]}}; // 10.0
    wire [7:0] v1848; shift_adder #(8, 2, 0, 0, 8, 0, 0) op_1848 (v1847[7:0], 2'b10, v1848[7:0]); // 10.0
    wire [4:0] v1849; assign v1849[4:0] = v1848[6:2]; // 10.0
    wire [8:0] v1850; shift_adder #(7, 8, 1, 1, 9, 0, 0) op_1850 (v1571[6:0], v1653[7:0], v1850[8:0]); // 10.0
    wire [8:0] v1851; shift_adder #(9, 2, 1, 0, 9, 0, 1) op_1851 (v1850[8:0], 2'b10, v1851[8:0]); // 10.0
    wire [7:0] v1852; assign v1852[7:0] = v1851[7:0] & {8{~v1851[8]}}; // 10.0
    wire [7:0] v1853; shift_adder #(8, 1, 0, 0, 8, 0, 0) op_1853 (v1852[7:0], 1'b1, v1853[7:0]); // 10.0
    wire [5:0] v1854; assign v1854[5:0] = v1853[6:1]; // 10.0
    wire [8:0] v1855; shift_adder #(8, 7, 1, 1, 9, 0, 0) op_1855 (v1573[7:0], v1654[6:0], v1855[8:0]); // 10.0
    wire [9:0] v1856; shift_adder #(9, 3, 1, 0, 10, -2, 1) op_1856 (v1855[8:0], 3'b101, v1856[9:0]); // 10.0
    wire [8:0] v1857; assign v1857[8:0] = v1856[8:0] & {9{~v1856[9]}}; // 10.0
    wire [8:0] v1858; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1858 (v1857[8:0], 3'b100, v1858[8:0]); // 10.0
    wire [5:0] v1859; assign v1859[5:0] = v1858[8:3]; // 10.0
    wire [9:0] v1860; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_1860 (v1655[7:0], v1656[7:0], v1860[9:0]); // 10.0
    wire [9:0] v1861; shift_adder #(10, 4, 1, 0, 10, -1, 0) op_1861 (v1860[9:0], 4'b1011, v1861[9:0]); // 10.0
    wire [8:0] v1862; assign v1862[8:0] = v1861[8:0] & {9{~v1861[9]}}; // 10.0
    wire [8:0] v1863; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1863 (v1862[8:0], 3'b100, v1863[8:0]); // 10.0
    wire [4:0] v1864; assign v1864[4:0] = v1863[7:3]; // 10.0
    wire [8:0] v1865; shift_adder #(8, 7, 1, 1, 9, 1, 0) op_1865 (v1577[7:0], v1657[6:0], v1865[8:0]); // 10.0
    wire [9:0] v1866; shift_adder #(9, 4, 1, 0, 10, -1, 1) op_1866 (v1865[8:0], 4'b1001, v1866[9:0]); // 10.0
    wire [8:0] v1867; assign v1867[8:0] = v1866[8:0] & {9{~v1866[9]}}; // 10.0
    wire [8:0] v1868; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1868 (v1867[8:0], 3'b100, v1868[8:0]); // 10.0
    wire [4:0] v1869; assign v1869[4:0] = v1868[7:3]; // 10.0
    wire [5:0] v1870; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_1870 (v1667[4:0], v1672[4:0], v1870[5:0]); // 10.0
    wire [6:0] v1871; shift_adder #(5, 5, 1, 1, 7, -1, 1) op_1871 (v1677[4:0], v1682[4:0], v1871[6:0]); // 10.0
    wire [9:0] v1872; shift_adder #(9, 7, 1, 1, 10, 1, 0) op_1872 (v1683[8:0], v1684[6:0], v1872[9:0]); // 10.0
    wire [9:0] v1873; shift_adder #(10, 4, 1, 0, 10, -1, 0) op_1873 (v1872[9:0], 4'b1011, v1873[9:0]); // 10.0
    wire [8:0] v1874; assign v1874[8:0] = v1873[8:0] & {9{~v1873[9]}}; // 10.0
    wire [8:0] v1875; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1875 (v1874[8:0], 3'b100, v1875[8:0]); // 10.0
    wire [4:0] v1876; assign v1876[4:0] = v1875[7:3]; // 10.0
    wire [9:0] v1877; shift_adder #(9, 8, 1, 1, 10, 1, 0) op_1877 (v1588[8:0], v1685[7:0], v1877[9:0]); // 10.0
    wire [9:0] v1878; shift_adder #(10, 3, 1, 0, 10, 0, 1) op_1878 (v1877[9:0], 3'b100, v1878[9:0]); // 10.0
    wire [8:0] v1879; assign v1879[8:0] = v1878[8:0] & {9{~v1878[9]}}; // 10.0
    wire [8:0] v1880; shift_adder #(9, 2, 0, 0, 9, 0, 0) op_1880 (v1879[8:0], 2'b10, v1880[8:0]); // 10.0
    wire [4:0] v1881; assign v1881[4:0] = v1880[6:2]; // 10.0
    wire [8:0] v1882; shift_adder #(7, 9, 1, 1, 9, -1, 0) op_1882 (v1590[6:0], v1686[8:0], v1882[8:0]); // 10.0
    wire [9:0] v1883; shift_adder #(9, 3, 1, 0, 10, -1, 1) op_1883 (v1882[8:0], 3'b101, v1883[9:0]); // 10.0
    wire [8:0] v1884; assign v1884[8:0] = v1883[8:0] & {9{~v1883[9]}}; // 10.0
    wire [8:0] v1885; shift_adder #(9, 3, 0, 0, 9, 0, 0) op_1885 (v1884[8:0], 3'b100, v1885[8:0]); // 10.0
    wire [4:0] v1886; assign v1886[4:0] = v1885[7:3]; // 10.0
    wire [8:0] v1887; shift_adder #(9, 7, 1, 1, 9, 1, 1) op_1887 (v1687[8:0], v1590[6:0], v1887[8:0]); // 10.0
    wire [8:0] v1888; shift_adder #(9, 3, 1, 0, 9, 0, 0) op_1888 (v1887[8:0], 3'b100, v1888[8:0]); // 10.0
    wire [7:0] v1889; assign v1889[7:0] = v1888[7:0] & {8{~v1888[8]}}; // 10.0
    wire [7:0] v1890; shift_adder #(8, 2, 0, 0, 8, 0, 0) op_1890 (v1889[7:0], 2'b10, v1890[7:0]); // 10.0
    wire [4:0] v1891; assign v1891[4:0] = v1890[6:2]; // 10.0
    wire [5:0] v1892; shift_adder #(4, 5, 1, 1, 6, -1, 0) op_1892 (v1597[3:0], v1692[4:0], v1892[5:0]); // 10.0
    wire [5:0] v1893; shift_adder #(5, 5, 1, 1, 6, 0, 0) op_1893 (v1697[4:0], v1610[4:0], v1893[5:0]); // 10.0
    wire [6:0] v1894; shift_adder #(4, 4, 1, 1, 7, -2, 1) op_1894 (v1630[3:0], v1702[3:0], v1894[6:0]); // 10.0
    wire [5:0] v1895; shift_adder #(5, 4, 1, 1, 6, 1, 0) op_1895 (v1707[4:0], v1630[3:0], v1895[5:0]); // 10.0
    wire [8:0] v1896; shift_adder #(7, 8, 1, 1, 9, 0, 0) op_1896 (v1603[6:0], v1708[7:0], v1896[8:0]); // 10.0
    wire [8:0] v1897; shift_adder #(9, 2, 1, 0, 9, 0, 1) op_1897 (v1896[8:0], 2'b10, v1897[8:0]); // 10.0
    wire [7:0] v1898; assign v1898[7:0] = v1897[7:0] & {8{~v1897[8]}}; // 10.0
    wire [7:0] v1899; shift_adder #(8, 1, 0, 0, 8, 0, 0) op_1899 (v1898[7:0], 1'b1, v1899[7:0]); // 10.0
    wire [5:0] v1900; assign v1900[5:0] = v1899[6:1]; // 10.0
    wire [6:0] v1901; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_1901 (v1667[4:0], v1672[4:0], v1901[6:0]); // 10.0
    wire [7:0] v1902; shift_adder #(5, 5, 1, 1, 8, -2, 1) op_1902 (v1682[4:0], v1682[4:0], v1902[7:0]); // 10.0
    wire [4:0] v1903; shift_adder #(4, 4, 1, 1, 5, 0, 0) op_1903 (v1630[3:0], v1702[3:0], v1903[4:0]); // 10.0
    wire [4:0] v1904; shift_adder #(4, 4, 1, 1, 5, 0, 1) op_1904 (v1625[3:0], v1597[3:0], v1904[4:0]); // 10.0
    wire [6:0] v1905; shift_adder #(5, 5, 1, 1, 7, 1, 0) op_1905 (v1692[4:0], v1610[4:0], v1905[6:0]); // 10.0
    wire [8:0] v1906; shift_adder #(5, 5, 1, 1, 9, -3, 0) op_1906 (v1707[4:0], v1697[4:0], v1906[8:0]); // 10.0

    // verilator lint_on UNUSEDSIGNAL

    assign model_out[4:0] = v1713[4:0];
    assign model_out[9:5] = v1610[4:0];
    assign model_out[15:10] = v1718[5:0];
    assign model_out[20:16] = v1723[4:0];
    assign model_out[25:21] = v1728[4:0];
    assign model_out[29:26] = v1733[3:0];
    assign model_out[34:30] = v1738[4:0];
    assign model_out[39:35] = v1743[4:0];
    assign model_out[44:40] = v1748[4:0];
    assign model_out[49:45] = v1753[4:0];
    assign model_out[54:50] = v1758[4:0];
    assign model_out[60:55] = v1759[5:0];
    assign model_out[65:61] = v1764[4:0];
    assign model_out[70:66] = v1769[4:0];
    assign model_out[76:71] = v1774[5:0];
    assign model_out[82:77] = v1779[5:0];
    assign model_out[87:83] = v1784[4:0];
    assign model_out[93:88] = v1789[5:0];
    assign model_out[98:94] = v1799[4:0];
    assign model_out[103:99] = v1804[4:0];
    assign model_out[108:104] = v1809[4:0];
    assign model_out[113:109] = v1814[4:0];
    assign model_out[119:114] = v1819[5:0];
    assign model_out[125:120] = v1824[5:0];
    assign model_out[130:126] = v1829[4:0];
    assign model_out[135:131] = v1834[4:0];
    assign model_out[140:136] = v1839[4:0];
    assign model_out[145:141] = v1844[4:0];
    assign model_out[150:146] = v1849[4:0];
    assign model_out[156:151] = v1854[5:0];
    assign model_out[162:157] = v1859[5:0];
    assign model_out[167:163] = v1864[4:0];
    assign model_out[172:168] = v1869[4:0];
    assign model_out[175:173] = v1662[2:0];
    assign model_out[181:176] = v1870[5:0];
    assign model_out[188:182] = v1871[6:0];
    assign model_out[193:189] = v1876[4:0];
    assign model_out[198:194] = v1881[4:0];
    assign model_out[203:199] = v1886[4:0];
    assign model_out[208:204] = v1891[4:0];
    assign model_out[214:209] = v1892[5:0];
    assign model_out[220:215] = v1893[5:0];
    assign model_out[227:221] = v1894[6:0];
    assign model_out[233:228] = v1895[5:0];
    assign model_out[240:234] = v1901[6:0];
    assign model_out[248:241] = v1902[7:0];
    assign model_out[254:249] = v1794[5:0];
    assign model_out[260:255] = v1900[5:0];
    assign model_out[265:261] = v1904[4:0];
    assign model_out[272:266] = v1905[6:0];
    assign model_out[281:273] = v1906[8:0];
    assign model_out[286:282] = v1903[4:0];

    endmodule
