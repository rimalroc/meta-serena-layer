`timescale 1 ns / 1 ps

module vmodel_stage0 (
    input [59:0] model_inp,
    output [69:0] model_out
);

    // verilator lint_off UNUSEDSIGNAL
    // Explicit quantization operation will drop bits if exists

    wire [0:0] v0; assign v0[0:0] = model_inp[0:0]; // 0.0
    wire [0:0] v1; assign v1[0:0] = model_inp[1:1]; // 0.0
    wire [0:0] v2; assign v2[0:0] = model_inp[2:2]; // 0.0
    wire [0:0] v3; assign v3[0:0] = model_inp[3:3]; // 0.0
    wire [0:0] v4; assign v4[0:0] = model_inp[4:4]; // 0.0
    wire [0:0] v5; assign v5[0:0] = model_inp[5:5]; // 0.0
    wire [0:0] v6; assign v6[0:0] = model_inp[6:6]; // 0.0
    wire [0:0] v7; assign v7[0:0] = model_inp[7:7]; // 0.0
    wire [0:0] v8; assign v8[0:0] = model_inp[8:8]; // 0.0
    wire [0:0] v9; assign v9[0:0] = model_inp[9:9]; // 0.0
    wire [0:0] v10; assign v10[0:0] = model_inp[10:10]; // 0.0
    wire [0:0] v11; assign v11[0:0] = model_inp[11:11]; // 0.0
    wire [0:0] v12; assign v12[0:0] = model_inp[12:12]; // 0.0
    wire [0:0] v13; assign v13[0:0] = model_inp[13:13]; // 0.0
    wire [0:0] v14; assign v14[0:0] = model_inp[14:14]; // 0.0
    wire [0:0] v15; assign v15[0:0] = model_inp[15:15]; // 0.0
    wire [0:0] v16; assign v16[0:0] = model_inp[16:16]; // 0.0
    wire [0:0] v17; assign v17[0:0] = model_inp[17:17]; // 0.0
    wire [0:0] v18; assign v18[0:0] = model_inp[18:18]; // 0.0
    wire [0:0] v19; assign v19[0:0] = model_inp[19:19]; // 0.0
    wire [0:0] v20; assign v20[0:0] = model_inp[20:20]; // 0.0
    wire [0:0] v21; assign v21[0:0] = model_inp[21:21]; // 0.0
    wire [0:0] v22; assign v22[0:0] = model_inp[22:22]; // 0.0
    wire [0:0] v23; assign v23[0:0] = model_inp[23:23]; // 0.0
    wire [0:0] v24; assign v24[0:0] = model_inp[24:24]; // 0.0
    wire [0:0] v25; assign v25[0:0] = model_inp[25:25]; // 0.0
    wire [0:0] v26; assign v26[0:0] = model_inp[26:26]; // 0.0
    wire [0:0] v27; assign v27[0:0] = model_inp[27:27]; // 0.0
    wire [0:0] v28; assign v28[0:0] = model_inp[28:28]; // 0.0
    wire [0:0] v29; assign v29[0:0] = model_inp[29:29]; // 0.0
    wire [0:0] v30; assign v30[0:0] = model_inp[30:30]; // 0.0
    wire [0:0] v31; assign v31[0:0] = model_inp[31:31]; // 0.0
    wire [0:0] v32; assign v32[0:0] = model_inp[32:32]; // 0.0
    wire [0:0] v33; assign v33[0:0] = model_inp[33:33]; // 0.0
    wire [0:0] v34; assign v34[0:0] = model_inp[34:34]; // 0.0
    wire [0:0] v35; assign v35[0:0] = model_inp[35:35]; // 0.0
    wire [0:0] v36; assign v36[0:0] = model_inp[36:36]; // 0.0
    wire [0:0] v37; assign v37[0:0] = model_inp[37:37]; // 0.0
    wire [0:0] v38; assign v38[0:0] = model_inp[38:38]; // 0.0
    wire [0:0] v39; assign v39[0:0] = model_inp[39:39]; // 0.0
    wire [0:0] v40; assign v40[0:0] = model_inp[40:40]; // 0.0
    wire [0:0] v41; assign v41[0:0] = model_inp[41:41]; // 0.0
    wire [0:0] v42; assign v42[0:0] = model_inp[42:42]; // 0.0
    wire [0:0] v43; assign v43[0:0] = model_inp[43:43]; // 0.0
    wire [0:0] v44; assign v44[0:0] = model_inp[44:44]; // 0.0
    wire [0:0] v45; assign v45[0:0] = model_inp[45:45]; // 0.0
    wire [0:0] v46; assign v46[0:0] = model_inp[46:46]; // 0.0
    wire [0:0] v47; assign v47[0:0] = model_inp[47:47]; // 0.0
    wire [0:0] v48; assign v48[0:0] = model_inp[48:48]; // 0.0
    wire [0:0] v49; assign v49[0:0] = model_inp[49:49]; // 0.0
    wire [0:0] v50; assign v50[0:0] = model_inp[50:50]; // 0.0
    wire [0:0] v51; assign v51[0:0] = model_inp[51:51]; // 0.0
    wire [0:0] v52; assign v52[0:0] = model_inp[52:52]; // 0.0
    wire [0:0] v53; assign v53[0:0] = model_inp[53:53]; // 0.0
    wire [0:0] v54; assign v54[0:0] = model_inp[54:54]; // 0.0
    wire [0:0] v55; assign v55[0:0] = model_inp[55:55]; // 0.0
    wire [0:0] v56; assign v56[0:0] = model_inp[56:56]; // 0.0
    wire [0:0] v57; assign v57[0:0] = model_inp[57:57]; // 0.0
    wire [0:0] v58; assign v58[0:0] = model_inp[58:58]; // 0.0
    wire [0:0] v59; assign v59[0:0] = model_inp[59:59]; // 0.0
    wire [0:0] v60; assign v60[0:0] = v0[0:0]; // 0.0
    wire [0:0] v61; assign v61[0:0] = v1[0:0]; // 0.0
    wire [0:0] v62; assign v62[0:0] = v2[0:0]; // 0.0
    wire [0:0] v63; assign v63[0:0] = v27[0:0]; // 0.0
    wire [0:0] v64; assign v64[0:0] = v28[0:0]; // 0.0
    wire [0:0] v65; assign v65[0:0] = v29[0:0]; // 0.0
    wire [0:0] v66; assign v66[0:0] = v33[0:0]; // 0.0
    wire [0:0] v67; assign v67[0:0] = v34[0:0]; // 0.0
    wire [0:0] v68; assign v68[0:0] = v35[0:0]; // 0.0
    wire [0:0] v69; assign v69[0:0] = v39[0:0]; // 0.0
    wire [0:0] v70; assign v70[0:0] = v40[0:0]; // 0.0
    wire [0:0] v71; assign v71[0:0] = v41[0:0]; // 0.0
    wire [0:0] v72; assign v72[0:0] = v45[0:0]; // 0.0
    wire [0:0] v73; assign v73[0:0] = v46[0:0]; // 0.0
    wire [0:0] v74; assign v74[0:0] = v47[0:0]; // 0.0
    wire [0:0] v75; assign v75[0:0] = v51[0:0]; // 0.0
    wire [0:0] v76; assign v76[0:0] = v52[0:0]; // 0.0
    wire [0:0] v77; assign v77[0:0] = v53[0:0]; // 0.0
    wire [0:0] v78; assign v78[0:0] = v57[0:0]; // 0.0
    wire [0:0] v79; assign v79[0:0] = v58[0:0]; // 0.0
    wire [0:0] v80; assign v80[0:0] = v59[0:0]; // 0.0
    wire [0:0] v81; assign v81[0:0] = v3[0:0]; // 0.0
    wire [0:0] v82; assign v82[0:0] = v4[0:0]; // 0.0
    wire [0:0] v83; assign v83[0:0] = v5[0:0]; // 0.0
    wire [0:0] v84; assign v84[0:0] = v9[0:0]; // 0.0
    wire [0:0] v85; assign v85[0:0] = v10[0:0]; // 0.0
    wire [0:0] v86; assign v86[0:0] = v11[0:0]; // 0.0
    wire [0:0] v87; assign v87[0:0] = v15[0:0]; // 0.0
    wire [0:0] v88; assign v88[0:0] = v16[0:0]; // 0.0
    wire [0:0] v89; assign v89[0:0] = v17[0:0]; // 0.0
    wire [0:0] v90; assign v90[0:0] = v21[0:0]; // 0.0
    wire [0:0] v91; assign v91[0:0] = v22[0:0]; // 0.0
    wire [0:0] v92; assign v92[0:0] = v23[0:0]; // 0.0
    wire [0:0] v93; assign v93[0:0] = v6[0:0]; // 0.0
    wire [0:0] v94; assign v94[0:0] = v7[0:0]; // 0.0
    wire [0:0] v95; assign v95[0:0] = v8[0:0]; // 0.0
    wire [0:0] v96; assign v96[0:0] = v12[0:0]; // 0.0
    wire [0:0] v97; assign v97[0:0] = v13[0:0]; // 0.0
    wire [0:0] v98; assign v98[0:0] = v14[0:0]; // 0.0
    wire [0:0] v99; assign v99[0:0] = v18[0:0]; // 0.0
    wire [0:0] v100; assign v100[0:0] = v19[0:0]; // 0.0
    wire [0:0] v101; assign v101[0:0] = v20[0:0]; // 0.0
    wire [0:0] v102; assign v102[0:0] = v24[0:0]; // 0.0
    wire [0:0] v103; assign v103[0:0] = v25[0:0]; // 0.0
    wire [0:0] v104; assign v104[0:0] = v26[0:0]; // 0.0
    wire [0:0] v105; assign v105[0:0] = v30[0:0]; // 0.0
    wire [0:0] v106; assign v106[0:0] = v31[0:0]; // 0.0
    wire [0:0] v107; assign v107[0:0] = v32[0:0]; // 0.0
    wire [0:0] v108; assign v108[0:0] = v36[0:0]; // 0.0
    wire [0:0] v109; assign v109[0:0] = v37[0:0]; // 0.0
    wire [0:0] v110; assign v110[0:0] = v38[0:0]; // 0.0
    wire [0:0] v111; assign v111[0:0] = v42[0:0]; // 0.0
    wire [0:0] v112; assign v112[0:0] = v43[0:0]; // 0.0
    wire [0:0] v113; assign v113[0:0] = v44[0:0]; // 0.0
    wire [0:0] v114; assign v114[0:0] = v48[0:0]; // 0.0
    wire [0:0] v115; assign v115[0:0] = v49[0:0]; // 0.0
    wire [0:0] v116; assign v116[0:0] = v50[0:0]; // 0.0
    wire [0:0] v117; assign v117[0:0] = v54[0:0]; // 0.0
    wire [0:0] v118; assign v118[0:0] = v55[0:0]; // 0.0
    wire [0:0] v119; assign v119[0:0] = v56[0:0]; // 0.0
    wire [1:0] v120; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_120 (v60[0:0], v61[0:0], v120[1:0]); // 1.0
    wire [1:0] v121; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_121 (v63[0:0], v64[0:0], v121[1:0]); // 1.0
    wire [1:0] v122; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_122 (v66[0:0], v67[0:0], v122[1:0]); // 1.0
    wire [1:0] v123; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_123 (v69[0:0], v70[0:0], v123[1:0]); // 1.0
    wire [1:0] v124; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_124 (v72[0:0], v73[0:0], v124[1:0]); // 1.0
    wire [1:0] v125; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_125 (v75[0:0], v76[0:0], v125[1:0]); // 1.0
    wire [1:0] v126; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_126 (v78[0:0], v79[0:0], v126[1:0]); // 1.0
    wire [1:0] v127; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_127 (v81[0:0], v82[0:0], v127[1:0]); // 1.0
    wire [1:0] v128; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_128 (v84[0:0], v85[0:0], v128[1:0]); // 1.0
    wire [1:0] v129; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_129 (v87[0:0], v88[0:0], v129[1:0]); // 1.0
    wire [1:0] v130; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_130 (v90[0:0], v91[0:0], v130[1:0]); // 1.0
    wire [1:0] v131; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_131 (v93[0:0], v94[0:0], v131[1:0]); // 1.0
    wire [1:0] v132; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_132 (v96[0:0], v97[0:0], v132[1:0]); // 1.0
    wire [1:0] v133; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_133 (v99[0:0], v100[0:0], v133[1:0]); // 1.0
    wire [1:0] v134; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_134 (v102[0:0], v103[0:0], v134[1:0]); // 1.0
    wire [1:0] v135; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_135 (v105[0:0], v106[0:0], v135[1:0]); // 1.0
    wire [1:0] v136; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_136 (v108[0:0], v109[0:0], v136[1:0]); // 1.0
    wire [1:0] v137; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_137 (v111[0:0], v112[0:0], v137[1:0]); // 1.0
    wire [1:0] v138; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_138 (v114[0:0], v115[0:0], v138[1:0]); // 1.0
    wire [1:0] v139; shift_adder #(1, 1, 0, 0, 2, 0, 0) op_139 (v117[0:0], v118[0:0], v139[1:0]); // 1.0
    wire [1:0] v140; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_140 (v120[1:0], v62[0:0], v140[1:0]); // 2.0
    wire [1:0] v141; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_141 (v121[1:0], v65[0:0], v141[1:0]); // 2.0
    wire [1:0] v142; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_142 (v122[1:0], v68[0:0], v142[1:0]); // 2.0
    wire [1:0] v143; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_143 (v123[1:0], v71[0:0], v143[1:0]); // 2.0
    wire [1:0] v144; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_144 (v124[1:0], v74[0:0], v144[1:0]); // 2.0
    wire [1:0] v145; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_145 (v125[1:0], v77[0:0], v145[1:0]); // 2.0
    wire [1:0] v146; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_146 (v126[1:0], v80[0:0], v146[1:0]); // 2.0
    wire [1:0] v147; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_147 (v127[1:0], v83[0:0], v147[1:0]); // 2.0
    wire [1:0] v148; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_148 (v128[1:0], v86[0:0], v148[1:0]); // 2.0
    wire [1:0] v149; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_149 (v129[1:0], v89[0:0], v149[1:0]); // 2.0
    wire [1:0] v150; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_150 (v130[1:0], v92[0:0], v150[1:0]); // 2.0
    wire [1:0] v151; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_151 (v131[1:0], v95[0:0], v151[1:0]); // 2.0
    wire [1:0] v152; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_152 (v132[1:0], v98[0:0], v152[1:0]); // 2.0
    wire [1:0] v153; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_153 (v133[1:0], v101[0:0], v153[1:0]); // 2.0
    wire [1:0] v154; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_154 (v134[1:0], v104[0:0], v154[1:0]); // 2.0
    wire [1:0] v155; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_155 (v135[1:0], v107[0:0], v155[1:0]); // 2.0
    wire [1:0] v156; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_156 (v136[1:0], v110[0:0], v156[1:0]); // 2.0
    wire [1:0] v157; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_157 (v137[1:0], v113[0:0], v157[1:0]); // 2.0
    wire [1:0] v158; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_158 (v138[1:0], v116[0:0], v158[1:0]); // 2.0
    wire [1:0] v159; shift_adder #(2, 1, 0, 0, 2, 0, 0) op_159 (v139[1:0], v119[0:0], v159[1:0]); // 2.0
    wire [3:0] v160; multiplier #(2, 2, 0, 0, 4) op_160 (v140[1:0], v141[1:0], v160[3:0]); // 4.0
    wire [3:0] v161; multiplier #(2, 2, 0, 0, 4) op_161 (v140[1:0], v142[1:0], v161[3:0]); // 4.0
    wire [3:0] v162; multiplier #(2, 2, 0, 0, 4) op_162 (v140[1:0], v143[1:0], v162[3:0]); // 4.0
    wire [3:0] v163; multiplier #(2, 2, 0, 0, 4) op_163 (v140[1:0], v144[1:0], v163[3:0]); // 4.0
    wire [3:0] v164; multiplier #(2, 2, 0, 0, 4) op_164 (v140[1:0], v145[1:0], v164[3:0]); // 4.0
    wire [3:0] v165; multiplier #(2, 2, 0, 0, 4) op_165 (v140[1:0], v146[1:0], v165[3:0]); // 4.0
    wire [3:0] v166; multiplier #(2, 2, 0, 0, 4) op_166 (v140[1:0], v147[1:0], v166[3:0]); // 4.0
    wire [3:0] v167; multiplier #(2, 2, 0, 0, 4) op_167 (v140[1:0], v148[1:0], v167[3:0]); // 4.0
    wire [3:0] v168; multiplier #(2, 2, 0, 0, 4) op_168 (v140[1:0], v149[1:0], v168[3:0]); // 4.0
    wire [3:0] v169; multiplier #(2, 2, 0, 0, 4) op_169 (v140[1:0], v150[1:0], v169[3:0]); // 4.0
    wire [3:0] v170; multiplier #(2, 2, 0, 0, 4) op_170 (v151[1:0], v141[1:0], v170[3:0]); // 4.0
    wire [3:0] v171; multiplier #(2, 2, 0, 0, 4) op_171 (v151[1:0], v142[1:0], v171[3:0]); // 4.0
    wire [3:0] v172; multiplier #(2, 2, 0, 0, 4) op_172 (v151[1:0], v143[1:0], v172[3:0]); // 4.0
    wire [3:0] v173; multiplier #(2, 2, 0, 0, 4) op_173 (v151[1:0], v144[1:0], v173[3:0]); // 4.0
    wire [3:0] v174; multiplier #(2, 2, 0, 0, 4) op_174 (v151[1:0], v145[1:0], v174[3:0]); // 4.0
    wire [3:0] v175; multiplier #(2, 2, 0, 0, 4) op_175 (v151[1:0], v146[1:0], v175[3:0]); // 4.0
    wire [3:0] v176; multiplier #(2, 2, 0, 0, 4) op_176 (v151[1:0], v147[1:0], v176[3:0]); // 4.0
    wire [3:0] v177; multiplier #(2, 2, 0, 0, 4) op_177 (v151[1:0], v148[1:0], v177[3:0]); // 4.0
    wire [3:0] v178; multiplier #(2, 2, 0, 0, 4) op_178 (v151[1:0], v149[1:0], v178[3:0]); // 4.0
    wire [3:0] v179; multiplier #(2, 2, 0, 0, 4) op_179 (v151[1:0], v150[1:0], v179[3:0]); // 4.0
    wire [3:0] v180; multiplier #(2, 2, 0, 0, 4) op_180 (v152[1:0], v141[1:0], v180[3:0]); // 4.0
    wire [3:0] v181; multiplier #(2, 2, 0, 0, 4) op_181 (v152[1:0], v142[1:0], v181[3:0]); // 4.0
    wire [3:0] v182; multiplier #(2, 2, 0, 0, 4) op_182 (v152[1:0], v143[1:0], v182[3:0]); // 4.0
    wire [3:0] v183; multiplier #(2, 2, 0, 0, 4) op_183 (v152[1:0], v144[1:0], v183[3:0]); // 4.0
    wire [3:0] v184; multiplier #(2, 2, 0, 0, 4) op_184 (v152[1:0], v145[1:0], v184[3:0]); // 4.0
    wire [3:0] v185; multiplier #(2, 2, 0, 0, 4) op_185 (v152[1:0], v146[1:0], v185[3:0]); // 4.0
    wire [3:0] v186; multiplier #(2, 2, 0, 0, 4) op_186 (v152[1:0], v147[1:0], v186[3:0]); // 4.0
    wire [3:0] v187; multiplier #(2, 2, 0, 0, 4) op_187 (v152[1:0], v148[1:0], v187[3:0]); // 4.0
    wire [3:0] v188; multiplier #(2, 2, 0, 0, 4) op_188 (v152[1:0], v149[1:0], v188[3:0]); // 4.0
    wire [3:0] v189; multiplier #(2, 2, 0, 0, 4) op_189 (v152[1:0], v150[1:0], v189[3:0]); // 4.0
    wire [3:0] v190; multiplier #(2, 2, 0, 0, 4) op_190 (v153[1:0], v141[1:0], v190[3:0]); // 4.0
    wire [3:0] v191; multiplier #(2, 2, 0, 0, 4) op_191 (v153[1:0], v142[1:0], v191[3:0]); // 4.0
    wire [3:0] v192; multiplier #(2, 2, 0, 0, 4) op_192 (v153[1:0], v143[1:0], v192[3:0]); // 4.0
    wire [3:0] v193; multiplier #(2, 2, 0, 0, 4) op_193 (v153[1:0], v144[1:0], v193[3:0]); // 4.0
    wire [3:0] v194; multiplier #(2, 2, 0, 0, 4) op_194 (v153[1:0], v145[1:0], v194[3:0]); // 4.0
    wire [3:0] v195; multiplier #(2, 2, 0, 0, 4) op_195 (v153[1:0], v146[1:0], v195[3:0]); // 4.0
    wire [3:0] v196; multiplier #(2, 2, 0, 0, 4) op_196 (v153[1:0], v147[1:0], v196[3:0]); // 4.0
    wire [3:0] v197; multiplier #(2, 2, 0, 0, 4) op_197 (v153[1:0], v148[1:0], v197[3:0]); // 4.0
    wire [3:0] v198; multiplier #(2, 2, 0, 0, 4) op_198 (v153[1:0], v149[1:0], v198[3:0]); // 4.0
    wire [3:0] v199; multiplier #(2, 2, 0, 0, 4) op_199 (v153[1:0], v150[1:0], v199[3:0]); // 4.0
    wire [3:0] v200; multiplier #(2, 2, 0, 0, 4) op_200 (v154[1:0], v141[1:0], v200[3:0]); // 4.0
    wire [3:0] v201; multiplier #(2, 2, 0, 0, 4) op_201 (v154[1:0], v142[1:0], v201[3:0]); // 4.0
    wire [3:0] v202; multiplier #(2, 2, 0, 0, 4) op_202 (v154[1:0], v143[1:0], v202[3:0]); // 4.0
    wire [3:0] v203; multiplier #(2, 2, 0, 0, 4) op_203 (v154[1:0], v144[1:0], v203[3:0]); // 4.0
    wire [3:0] v204; multiplier #(2, 2, 0, 0, 4) op_204 (v154[1:0], v145[1:0], v204[3:0]); // 4.0
    wire [3:0] v205; multiplier #(2, 2, 0, 0, 4) op_205 (v154[1:0], v146[1:0], v205[3:0]); // 4.0
    wire [3:0] v206; multiplier #(2, 2, 0, 0, 4) op_206 (v154[1:0], v147[1:0], v206[3:0]); // 4.0
    wire [3:0] v207; multiplier #(2, 2, 0, 0, 4) op_207 (v154[1:0], v148[1:0], v207[3:0]); // 4.0
    wire [3:0] v208; multiplier #(2, 2, 0, 0, 4) op_208 (v154[1:0], v149[1:0], v208[3:0]); // 4.0
    wire [3:0] v209; multiplier #(2, 2, 0, 0, 4) op_209 (v154[1:0], v150[1:0], v209[3:0]); // 4.0
    wire [3:0] v210; multiplier #(2, 2, 0, 0, 4) op_210 (v155[1:0], v141[1:0], v210[3:0]); // 4.0
    wire [3:0] v211; multiplier #(2, 2, 0, 0, 4) op_211 (v155[1:0], v142[1:0], v211[3:0]); // 4.0
    wire [3:0] v212; multiplier #(2, 2, 0, 0, 4) op_212 (v155[1:0], v143[1:0], v212[3:0]); // 4.0
    wire [3:0] v213; multiplier #(2, 2, 0, 0, 4) op_213 (v155[1:0], v144[1:0], v213[3:0]); // 4.0
    wire [3:0] v214; multiplier #(2, 2, 0, 0, 4) op_214 (v155[1:0], v145[1:0], v214[3:0]); // 4.0
    wire [3:0] v215; multiplier #(2, 2, 0, 0, 4) op_215 (v155[1:0], v146[1:0], v215[3:0]); // 4.0
    wire [3:0] v216; multiplier #(2, 2, 0, 0, 4) op_216 (v155[1:0], v147[1:0], v216[3:0]); // 4.0
    wire [3:0] v217; multiplier #(2, 2, 0, 0, 4) op_217 (v155[1:0], v148[1:0], v217[3:0]); // 4.0
    wire [3:0] v218; multiplier #(2, 2, 0, 0, 4) op_218 (v155[1:0], v149[1:0], v218[3:0]); // 4.0
    wire [3:0] v219; multiplier #(2, 2, 0, 0, 4) op_219 (v155[1:0], v150[1:0], v219[3:0]); // 4.0
    wire [3:0] v220; multiplier #(2, 2, 0, 0, 4) op_220 (v156[1:0], v141[1:0], v220[3:0]); // 4.0
    wire [3:0] v221; multiplier #(2, 2, 0, 0, 4) op_221 (v156[1:0], v142[1:0], v221[3:0]); // 4.0
    wire [3:0] v222; multiplier #(2, 2, 0, 0, 4) op_222 (v156[1:0], v143[1:0], v222[3:0]); // 4.0
    wire [3:0] v223; multiplier #(2, 2, 0, 0, 4) op_223 (v156[1:0], v144[1:0], v223[3:0]); // 4.0
    wire [3:0] v224; multiplier #(2, 2, 0, 0, 4) op_224 (v156[1:0], v145[1:0], v224[3:0]); // 4.0
    wire [3:0] v225; multiplier #(2, 2, 0, 0, 4) op_225 (v156[1:0], v146[1:0], v225[3:0]); // 4.0
    wire [3:0] v226; multiplier #(2, 2, 0, 0, 4) op_226 (v156[1:0], v147[1:0], v226[3:0]); // 4.0
    wire [3:0] v227; multiplier #(2, 2, 0, 0, 4) op_227 (v156[1:0], v148[1:0], v227[3:0]); // 4.0
    wire [3:0] v228; multiplier #(2, 2, 0, 0, 4) op_228 (v156[1:0], v149[1:0], v228[3:0]); // 4.0
    wire [3:0] v229; multiplier #(2, 2, 0, 0, 4) op_229 (v156[1:0], v150[1:0], v229[3:0]); // 4.0
    wire [3:0] v230; multiplier #(2, 2, 0, 0, 4) op_230 (v157[1:0], v141[1:0], v230[3:0]); // 4.0
    wire [3:0] v231; multiplier #(2, 2, 0, 0, 4) op_231 (v157[1:0], v142[1:0], v231[3:0]); // 4.0
    wire [3:0] v232; multiplier #(2, 2, 0, 0, 4) op_232 (v157[1:0], v143[1:0], v232[3:0]); // 4.0
    wire [3:0] v233; multiplier #(2, 2, 0, 0, 4) op_233 (v157[1:0], v144[1:0], v233[3:0]); // 4.0
    wire [3:0] v234; multiplier #(2, 2, 0, 0, 4) op_234 (v157[1:0], v145[1:0], v234[3:0]); // 4.0
    wire [3:0] v235; multiplier #(2, 2, 0, 0, 4) op_235 (v157[1:0], v146[1:0], v235[3:0]); // 4.0
    wire [3:0] v236; multiplier #(2, 2, 0, 0, 4) op_236 (v157[1:0], v147[1:0], v236[3:0]); // 4.0
    wire [3:0] v237; multiplier #(2, 2, 0, 0, 4) op_237 (v157[1:0], v148[1:0], v237[3:0]); // 4.0
    wire [3:0] v238; multiplier #(2, 2, 0, 0, 4) op_238 (v157[1:0], v149[1:0], v238[3:0]); // 4.0
    wire [3:0] v239; multiplier #(2, 2, 0, 0, 4) op_239 (v157[1:0], v150[1:0], v239[3:0]); // 4.0
    wire [3:0] v240; multiplier #(2, 2, 0, 0, 4) op_240 (v158[1:0], v141[1:0], v240[3:0]); // 4.0
    wire [3:0] v241; multiplier #(2, 2, 0, 0, 4) op_241 (v158[1:0], v142[1:0], v241[3:0]); // 4.0
    wire [3:0] v242; multiplier #(2, 2, 0, 0, 4) op_242 (v158[1:0], v143[1:0], v242[3:0]); // 4.0
    wire [3:0] v243; multiplier #(2, 2, 0, 0, 4) op_243 (v158[1:0], v144[1:0], v243[3:0]); // 4.0
    wire [3:0] v244; multiplier #(2, 2, 0, 0, 4) op_244 (v158[1:0], v145[1:0], v244[3:0]); // 4.0
    wire [3:0] v245; multiplier #(2, 2, 0, 0, 4) op_245 (v158[1:0], v146[1:0], v245[3:0]); // 4.0
    wire [3:0] v246; multiplier #(2, 2, 0, 0, 4) op_246 (v158[1:0], v147[1:0], v246[3:0]); // 4.0
    wire [3:0] v247; multiplier #(2, 2, 0, 0, 4) op_247 (v158[1:0], v148[1:0], v247[3:0]); // 4.0
    wire [3:0] v248; multiplier #(2, 2, 0, 0, 4) op_248 (v158[1:0], v149[1:0], v248[3:0]); // 4.0
    wire [3:0] v249; multiplier #(2, 2, 0, 0, 4) op_249 (v158[1:0], v150[1:0], v249[3:0]); // 4.0
    wire [3:0] v250; multiplier #(2, 2, 0, 0, 4) op_250 (v159[1:0], v141[1:0], v250[3:0]); // 4.0
    wire [3:0] v251; multiplier #(2, 2, 0, 0, 4) op_251 (v159[1:0], v142[1:0], v251[3:0]); // 4.0
    wire [3:0] v252; multiplier #(2, 2, 0, 0, 4) op_252 (v159[1:0], v143[1:0], v252[3:0]); // 4.0
    wire [3:0] v253; multiplier #(2, 2, 0, 0, 4) op_253 (v159[1:0], v144[1:0], v253[3:0]); // 4.0
    wire [3:0] v254; multiplier #(2, 2, 0, 0, 4) op_254 (v159[1:0], v145[1:0], v254[3:0]); // 4.0
    wire [3:0] v255; multiplier #(2, 2, 0, 0, 4) op_255 (v159[1:0], v146[1:0], v255[3:0]); // 4.0
    wire [3:0] v256; multiplier #(2, 2, 0, 0, 4) op_256 (v159[1:0], v147[1:0], v256[3:0]); // 4.0
    wire [3:0] v257; multiplier #(2, 2, 0, 0, 4) op_257 (v159[1:0], v148[1:0], v257[3:0]); // 4.0
    wire [3:0] v258; multiplier #(2, 2, 0, 0, 4) op_258 (v159[1:0], v149[1:0], v258[3:0]); // 4.0
    wire [3:0] v259; multiplier #(2, 2, 0, 0, 4) op_259 (v159[1:0], v150[1:0], v259[3:0]); // 4.0
    wire [4:0] v260; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_260 (v160[3:0], v161[3:0], v260[4:0]); // 5.0
    wire [4:0] v261; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_261 (v162[3:0], v163[3:0], v261[4:0]); // 5.0
    wire [4:0] v262; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_262 (v164[3:0], v165[3:0], v262[4:0]); // 5.0
    wire [4:0] v263; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_263 (v166[3:0], v167[3:0], v263[4:0]); // 5.0
    wire [4:0] v264; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_264 (v168[3:0], v169[3:0], v264[4:0]); // 5.0
    wire [4:0] v265; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_265 (v170[3:0], v171[3:0], v265[4:0]); // 5.0
    wire [4:0] v266; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_266 (v172[3:0], v173[3:0], v266[4:0]); // 5.0
    wire [4:0] v267; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_267 (v174[3:0], v175[3:0], v267[4:0]); // 5.0
    wire [4:0] v268; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_268 (v176[3:0], v177[3:0], v268[4:0]); // 5.0
    wire [4:0] v269; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_269 (v178[3:0], v179[3:0], v269[4:0]); // 5.0
    wire [4:0] v270; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_270 (v180[3:0], v181[3:0], v270[4:0]); // 5.0
    wire [4:0] v271; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_271 (v182[3:0], v183[3:0], v271[4:0]); // 5.0
    wire [4:0] v272; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_272 (v184[3:0], v185[3:0], v272[4:0]); // 5.0
    wire [4:0] v273; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_273 (v186[3:0], v187[3:0], v273[4:0]); // 5.0
    wire [4:0] v274; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_274 (v188[3:0], v189[3:0], v274[4:0]); // 5.0
    wire [4:0] v275; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_275 (v190[3:0], v191[3:0], v275[4:0]); // 5.0
    wire [4:0] v276; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_276 (v192[3:0], v193[3:0], v276[4:0]); // 5.0
    wire [4:0] v277; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_277 (v194[3:0], v195[3:0], v277[4:0]); // 5.0
    wire [4:0] v278; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_278 (v196[3:0], v197[3:0], v278[4:0]); // 5.0
    wire [4:0] v279; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_279 (v198[3:0], v199[3:0], v279[4:0]); // 5.0
    wire [4:0] v280; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_280 (v200[3:0], v201[3:0], v280[4:0]); // 5.0
    wire [4:0] v281; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_281 (v202[3:0], v203[3:0], v281[4:0]); // 5.0
    wire [4:0] v282; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_282 (v204[3:0], v205[3:0], v282[4:0]); // 5.0
    wire [4:0] v283; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_283 (v206[3:0], v207[3:0], v283[4:0]); // 5.0
    wire [4:0] v284; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_284 (v208[3:0], v209[3:0], v284[4:0]); // 5.0
    wire [4:0] v285; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_285 (v210[3:0], v211[3:0], v285[4:0]); // 5.0
    wire [4:0] v286; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_286 (v212[3:0], v213[3:0], v286[4:0]); // 5.0
    wire [4:0] v287; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_287 (v214[3:0], v215[3:0], v287[4:0]); // 5.0
    wire [4:0] v288; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_288 (v216[3:0], v217[3:0], v288[4:0]); // 5.0
    wire [4:0] v289; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_289 (v218[3:0], v219[3:0], v289[4:0]); // 5.0
    wire [4:0] v290; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_290 (v220[3:0], v221[3:0], v290[4:0]); // 5.0
    wire [4:0] v291; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_291 (v222[3:0], v223[3:0], v291[4:0]); // 5.0
    wire [4:0] v292; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_292 (v224[3:0], v225[3:0], v292[4:0]); // 5.0
    wire [4:0] v293; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_293 (v226[3:0], v227[3:0], v293[4:0]); // 5.0
    wire [4:0] v294; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_294 (v228[3:0], v229[3:0], v294[4:0]); // 5.0
    wire [4:0] v295; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_295 (v230[3:0], v231[3:0], v295[4:0]); // 5.0
    wire [4:0] v296; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_296 (v232[3:0], v233[3:0], v296[4:0]); // 5.0
    wire [4:0] v297; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_297 (v234[3:0], v235[3:0], v297[4:0]); // 5.0
    wire [4:0] v298; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_298 (v236[3:0], v237[3:0], v298[4:0]); // 5.0
    wire [4:0] v299; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_299 (v238[3:0], v239[3:0], v299[4:0]); // 5.0
    wire [4:0] v300; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_300 (v240[3:0], v241[3:0], v300[4:0]); // 5.0
    wire [4:0] v301; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_301 (v242[3:0], v243[3:0], v301[4:0]); // 5.0
    wire [4:0] v302; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_302 (v244[3:0], v245[3:0], v302[4:0]); // 5.0
    wire [4:0] v303; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_303 (v246[3:0], v247[3:0], v303[4:0]); // 5.0
    wire [4:0] v304; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_304 (v248[3:0], v249[3:0], v304[4:0]); // 5.0
    wire [4:0] v305; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_305 (v250[3:0], v251[3:0], v305[4:0]); // 5.0
    wire [4:0] v306; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_306 (v252[3:0], v253[3:0], v306[4:0]); // 5.0
    wire [4:0] v307; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_307 (v254[3:0], v255[3:0], v307[4:0]); // 5.0
    wire [4:0] v308; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_308 (v256[3:0], v257[3:0], v308[4:0]); // 5.0
    wire [4:0] v309; shift_adder #(4, 4, 0, 0, 5, 0, 0) op_309 (v258[3:0], v259[3:0], v309[4:0]); // 5.0
    wire [5:0] v310; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_310 (v260[4:0], v261[4:0], v310[5:0]); // 6.0
    wire [5:0] v311; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_311 (v263[4:0], v264[4:0], v311[5:0]); // 6.0
    wire [5:0] v312; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_312 (v265[4:0], v266[4:0], v312[5:0]); // 6.0
    wire [5:0] v313; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_313 (v268[4:0], v269[4:0], v313[5:0]); // 6.0
    wire [5:0] v314; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_314 (v270[4:0], v271[4:0], v314[5:0]); // 6.0
    wire [5:0] v315; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_315 (v273[4:0], v274[4:0], v315[5:0]); // 6.0
    wire [5:0] v316; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_316 (v275[4:0], v276[4:0], v316[5:0]); // 6.0
    wire [5:0] v317; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_317 (v278[4:0], v279[4:0], v317[5:0]); // 6.0
    wire [5:0] v318; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_318 (v280[4:0], v281[4:0], v318[5:0]); // 6.0
    wire [5:0] v319; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_319 (v283[4:0], v284[4:0], v319[5:0]); // 6.0
    wire [5:0] v320; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_320 (v285[4:0], v286[4:0], v320[5:0]); // 6.0
    wire [5:0] v321; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_321 (v288[4:0], v289[4:0], v321[5:0]); // 6.0
    wire [5:0] v322; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_322 (v290[4:0], v291[4:0], v322[5:0]); // 6.0
    wire [5:0] v323; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_323 (v293[4:0], v294[4:0], v323[5:0]); // 6.0
    wire [5:0] v324; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_324 (v295[4:0], v296[4:0], v324[5:0]); // 6.0
    wire [5:0] v325; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_325 (v298[4:0], v299[4:0], v325[5:0]); // 6.0
    wire [5:0] v326; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_326 (v300[4:0], v301[4:0], v326[5:0]); // 6.0
    wire [5:0] v327; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_327 (v303[4:0], v304[4:0], v327[5:0]); // 6.0
    wire [5:0] v328; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_328 (v305[4:0], v306[4:0], v328[5:0]); // 6.0
    wire [5:0] v329; shift_adder #(5, 5, 0, 0, 6, 0, 0) op_329 (v308[4:0], v309[4:0], v329[5:0]); // 6.0
    wire [5:0] v330; shift_adder #(5, 6, 0, 0, 6, 0, 0) op_330 (v262[4:0], v311[5:0], v330[5:0]); // 7.0
    wire [5:0] v331; shift_adder #(5, 6, 0, 0, 6, 0, 0) op_331 (v267[4:0], v313[5:0], v331[5:0]); // 7.0
    wire [5:0] v332; shift_adder #(5, 6, 0, 0, 6, 0, 0) op_332 (v272[4:0], v315[5:0], v332[5:0]); // 7.0
    wire [5:0] v333; shift_adder #(5, 6, 0, 0, 6, 0, 0) op_333 (v277[4:0], v317[5:0], v333[5:0]); // 7.0
    wire [5:0] v334; shift_adder #(5, 6, 0, 0, 6, 0, 0) op_334 (v282[4:0], v319[5:0], v334[5:0]); // 7.0
    wire [5:0] v335; shift_adder #(5, 6, 0, 0, 6, 0, 0) op_335 (v287[4:0], v321[5:0], v335[5:0]); // 7.0
    wire [5:0] v336; shift_adder #(5, 6, 0, 0, 6, 0, 0) op_336 (v292[4:0], v323[5:0], v336[5:0]); // 7.0
    wire [5:0] v337; shift_adder #(5, 6, 0, 0, 6, 0, 0) op_337 (v297[4:0], v325[5:0], v337[5:0]); // 7.0
    wire [5:0] v338; shift_adder #(5, 6, 0, 0, 6, 0, 0) op_338 (v302[4:0], v327[5:0], v338[5:0]); // 7.0
    wire [5:0] v339; shift_adder #(5, 6, 0, 0, 6, 0, 0) op_339 (v307[4:0], v329[5:0], v339[5:0]); // 7.0
    wire [6:0] v340; shift_adder #(6, 6, 0, 0, 7, 0, 0) op_340 (v310[5:0], v330[5:0], v340[6:0]); // 8.0
    wire [6:0] v341; shift_adder #(6, 6, 0, 0, 7, 0, 0) op_341 (v312[5:0], v331[5:0], v341[6:0]); // 8.0
    wire [6:0] v342; shift_adder #(6, 6, 0, 0, 7, 0, 0) op_342 (v314[5:0], v332[5:0], v342[6:0]); // 8.0
    wire [6:0] v343; shift_adder #(6, 6, 0, 0, 7, 0, 0) op_343 (v316[5:0], v333[5:0], v343[6:0]); // 8.0
    wire [6:0] v344; shift_adder #(6, 6, 0, 0, 7, 0, 0) op_344 (v318[5:0], v334[5:0], v344[6:0]); // 8.0
    wire [6:0] v345; shift_adder #(6, 6, 0, 0, 7, 0, 0) op_345 (v320[5:0], v335[5:0], v345[6:0]); // 8.0
    wire [6:0] v346; shift_adder #(6, 6, 0, 0, 7, 0, 0) op_346 (v322[5:0], v336[5:0], v346[6:0]); // 8.0
    wire [6:0] v347; shift_adder #(6, 6, 0, 0, 7, 0, 0) op_347 (v324[5:0], v337[5:0], v347[6:0]); // 8.0
    wire [6:0] v348; shift_adder #(6, 6, 0, 0, 7, 0, 0) op_348 (v326[5:0], v338[5:0], v348[6:0]); // 8.0
    wire [6:0] v349; shift_adder #(6, 6, 0, 0, 7, 0, 0) op_349 (v328[5:0], v339[5:0], v349[6:0]); // 8.0

    // verilator lint_on UNUSEDSIGNAL

    assign model_out[6:0] = v340[6:0];
    assign model_out[13:7] = v341[6:0];
    assign model_out[20:14] = v342[6:0];
    assign model_out[27:21] = v343[6:0];
    assign model_out[34:28] = v344[6:0];
    assign model_out[41:35] = v345[6:0];
    assign model_out[48:42] = v346[6:0];
    assign model_out[55:49] = v347[6:0];
    assign model_out[62:56] = v348[6:0];
    assign model_out[69:63] = v349[6:0];

    endmodule
